Vim�UnDo� oc?1�n�$s��p��M���q��P
��XxC�  _   int iter_k;   k   
     m      m  m  m    Z5�   " _�                            ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �                �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �                   �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �         !          �              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �         !    �         !    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �         "    �         "    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �          #    �         #    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �         $              rand logic espresso;5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �         $              rand logic espresso;5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             Z5	�     �          $              rand logic espresso;5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             Z5
     �         $              rand logic espresso;5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             Z5
     �         $              rand logic milk;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5
     �         $              rand logic chocolate;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5
     �          $              rand logic froth;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z5
>     �      "   %              �      !   $    5�_�                    !       ����                                                                                                                                                                                                                                                                                                                                                             Z5
E     �       "   &              rand logic5�_�                    !       ����                                                                                                                                                                                                                                                                                                                                                             Z5
E     �       "   &              rand logic[]5�_�                    !       ����                                                                                                                                                                                                                                                                                                                                                             Z5
G     �       "   &              rand logic[]5�_�                    !       ����                                                                                                                                                                                                                                                                                                                                                             Z5
I     �       "   &              rand logic[9:0]5�_�                    !   '    ����                                                                                                                                                                                                                                                                                                                                                             Z5
]     �   !   #   &    �   !   "   &    5�_�                    "       ����                                                                                                                                                                                                                                                                                                                                                             Z5
^     �   "   $   '    �   "   #   '    5�_�                    #       ����                                                                                                                                                                                                                                                                                                                                                             Z5
^     �   #   %   (    �   #   $   (    5�_�                    "       ����                                                                                                                                                                                                                                                                                                                                                             Z5
c     �   !   #   )      (        rand logic[9:0] espresso_addnum;5�_�                    "       ����                                                                                                                                                                                                                                                                                                                                                             Z5
d     �   !   #   )               rand logic[9:0] _addnum;5�_�                    "       ����                                                                                                                                                                                                                                                                                                                                                             Z5
f     �   !   #   )               rand logic[9:0] _addnum;5�_�                    #       ����                                                                                                                                                                                                                                                                                                                                                             Z5
i     �   "   $   )      (        rand logic[9:0] espresso_addnum;5�_�                    #       ����                                                                                                                                                                                                                                                                                                                                                             Z5
i     �   "   $   )               rand logic[9:0] _addnum;5�_�                    #       ����                                                                                                                                                                                                                                                                                                                                                             Z5
j     �   "   $   )               rand logic[9:0] _addnum;5�_�                    $       ����                                                                                                                                                                                                                                                                                                                                                             Z5
m     �   #   %   )      (        rand logic[9:0] espresso_addnum;5�_�                    $       ����                                                                                                                                                                                                                                                                                                                                                             Z5
m     �   #   %   )               rand logic[9:0] _addnum;5�_�                    $       ����                                                                                                                                                                                                                                                                                                                                                             Z5
n    �   #   %   )               rand logic[9:0] _addnum;5�_�                     %        ����                                                                                                                                                                                                                                                                                                                                                             Z5
�     �   $   %           5�_�      !               %        ����                                                                                                                                                                                                                                                                                                                                                             Z5
�     �   %   '   )              �   %   '   (    5�_�       "           !   &       ����                                                                                                                                                                                                                                                                                                                                                             Z5
�     �   %   )   )              constraint limit5�_�   !   #           "   (       ����                                                                                                                                                                                                                                                                                                                                                             Z5
�     �   '   )   +      	        }5�_�   "   $           #   '       ����                                                                                                                                                                                                                                                                                                                                                             Z5
�     �   &   (   +              5�_�   #   &           $   $   %    ����                                                                                                                                                                                                                                                                                                                            !          $   %          &    Z5     �   #   %   +      %        rand logic[9:0] froth_addnum;5�_�   $   '   %       &   '       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   '   ,   ,              �   '   )   +    5�_�   &   (           '   (        ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   '   )   /       5�_�   '   )           (   (       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   '   -   /                                 	        }�   (   )   /    5�_�   (   *           )   '       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   &   '                       espresso_addnum > 0;5�_�   )   +           *   '       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   &   (   .                  espresso_addnum;5�_�   *   ,           +   (       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   '   )   .                  milk_addnum;5�_�   +   -           ,   )       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   (   *   .                  chocolate_addnum5�_�   ,   .           -   *       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5!    �   )   +   .                  froth_addnum;   5�_�   -   /           .   ,       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5+     �   ,   0   /       �   ,   .   .    5�_�   .   0           /   /       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5>     �   /   1   1    5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5B     �         2      class supply_cl;5�_�   0   2           1   /       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5r     �   /   2   3          �   /   1   2    5�_�   1   3           2   /       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5u     �   /   1   5          �   /   1   4    5�_�   2   4           3   0       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   0   2   6              �   0   2   5    5�_�   3   5           4   1       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   0   1                      this.srandomdd5�_�   4   6           5   0        ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   0   2   6              �   0   2   5    5�_�   5   7           6   1       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   0   4   6              constraint5�_�   6   8           7   3       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   2   4   8      	        }5�_�   7   9           8   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   1   3   8              5�_�   8   :           9   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   1   3   8                  flavo5�_�   9   ;           :   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   1   3   8                  flavor_in inside 5�_�   :   <           ;   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   1   3   8                  flavor_in inside {}5�_�   ;   =           <   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   1   3   8                  flavor_in inside {}5�_�   <   >           =   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   1   3   8                  flavor_in inside {}5�_�   =   ?           >   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5�     �   1   3   8                  flavor_in inside {}5�_�   >   @           ?   0       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   0   2   9              �   0   2   8    5�_�   ?   A           @   1       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   0   2   9              function new5�_�   @   B           A   1       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   0   2   9              function new()5�_�   A   C           B   1       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   0   2   9              function new()5�_�   B   D           C   1       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   0   4   9              function new(int seed)5�_�   C   E           D   2        ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   1   3   ;       5�_�   D   F           E   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   1   3   ;                      this.srandom5�_�   E   G           F   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   1   3   ;                      this.srandom()5�_�   F   H           G   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   1   3   ;                      this.srandom()5�_�   G   I           H   2   "    ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5"    �   1   3   ;      "                this.srandom(seed)5�_�   H   J           I   4       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5(     �   3   5   ;              constraint{5�_�   I   K           J   7        ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5-     �   6   7           5�_�   J   L           K   0       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z50     �   0   2   :    5�_�   K   M           L   4       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z51     �   4   6   <              �   4   6   ;    5�_�   L   N           M   2       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z54     �   1   3   <              function new(int seed);5�_�   M   O           N   %        ����                                                                                                                                                                                                                                                                                                                            2   %       4          V   %    Z5E     �   %   )   <    �   %   &   <    5�_�   N   P           O   (       ����                                                                                                                                                                                                                                                                                                                            5   %       7          V   %    Z5F    �   (   *   ?    5�_�   O   Q           P   >        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5q     �   >   m   @    �   >   ?   @    5�_�   P   R           Q   @        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5x     �   ?   @              randc flavor flavor_in;5�_�   Q   S           R   @       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5y     �   ?   @              function new(int seed);5�_�   R   T           S   @       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5y     �   ?   @                      this.srandom(seed);5�_�   S   U           T   @       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5z     �   ?   @              endfunction 5�_�   T   V           U   @       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5z     �   ?   @              constraint limit 5�_�   U   W           V   @       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5z     �   ?   @              {5�_�   V   X           W   @       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5z     �   ?   @          6        !(flavor_in inside{no_coffee, 'd5, 'd6, 'd7});5�_�   W   Y           X   @       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5z     �   ?   @              }5�_�   X   Z           Y   @        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5{     �   ?   @          endclass5�_�   Y   [           Z   ?        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5{     �   >   ?          class select_flavor;5�_�   Z   \           [   3        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5}     �   3   5   d    �   3   4   d    5�_�   [   ]           \   3        ����                                                                                                                                                                                                                                                                                                                            7   %       9          V   %    Z5~     �   2   3          class flavor_rand;5�_�   \   ^           ]   ;   5    ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   :   <   d      5            flavor_in inside {latte,cappuccino,mocha}5�_�   ]   _           ^   ;   5    ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   :   <   d      5            flavor_in inside {latte,cappuccino,mocha}5�_�   ^   `           _   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              rand logic[2:0] espresso;5�_�   _   a           `   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              rand logic[2:0] milk;5�_�   `   b           a   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              rand logic[2:0] chocolate;5�_�   a   c           b   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              rand logic[2:0] froth;5�_�   b   d           c   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              function new(int seed);5�_�   c   e           d   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L                      this.srandom(seed);5�_�   d   f           e   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              endfunction 5�_�   e   g           f   K       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   M   ^          �   K   M   ]    5�_�   f   h           g   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              j5�_�   g   i           h   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              constraint limit 5�_�   h   j           i   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              {5�_�   i   k           j   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L          0        espresso + milk + chocolate + froth > 0;5�_�   j   l           k   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              }5�_�   k   m           l   K        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   M   Z          �   K   M   Y    5�_�   l   n           m   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   M   Z          function getratio5�_�   m   o           n   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   M   Z          function getratio()5�_�   n   p           o   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   L   O   [              �   L   N   Z    5�_�   o   q           p   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   L   N   ]              �   L   N   \    5�_�   p   r           q   N        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   M   N           5�_�   q   s           r   K       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   M   ]          �   K   M   \    5�_�   r   t           s   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5      �   K   M   ]          5�_�   s   u           t   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5     �   K   L              5�_�   t   v           u   K       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z50     �   K   M   \    5�_�   u   w           v   L        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z52     �   K   M   ]       5�_�   v   x           w   L   
    ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z51     �   K   M   ]      
    logic 5�_�   w   y           x   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z51     �   K   M   ]          logic []5�_�   x   z           y   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z54     �   K   M   ]          logic []5�_�   y   {           z   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z55     �   K   M   ]          logic [3:0]5�_�   z   |           {   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z57     �   K   M   ]          logic [2:0]5�_�   {   }           |   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z57     �   K   M   ]          logic [2:0]5�_�   |   ~           }   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5B     �   L   N   ]    �   L   M   ]    5�_�   }              ~   M       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5D     �   L   N   ^          logic [2:0] x_value;5�_�   ~   �              M       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5M     �   M   P   _          �   M   O   ^    5�_�      �           �   N        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5O     �   M   O   `       5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5T     �   M   O   `          function new5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5T     �   M   O   `          function new()5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5U     �   N   Q   a              �   N   P   `    5�_�   �   �           �   O        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5Z     �   N   P   b       5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5c     �   O   Q   b    �   O   P   b    5�_�   �   �           �   P       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5e     �   O   Q   c              this.x_value = 0;5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5i     �   S   T                  return5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5j     �   S   U   c              �   S   U   b    5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5w     �   S   U   c              this.y_value = 5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5w     �   S   U   c              this.y_value = ()5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5x     �   S   U   c              this.y_value = ()5�_�   �   �           �   T   *    ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   U   c      *        this.y_value = (this.y_value == 7)5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   U   c      @        this.y_value = (this.y_value == 7) ? 0 : this.y_value++;5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   U   c      <        .y_value = (this.y_value == 7) ? 0 : this.y_value++;5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   U   c      ;        y_value = (this.y_value == 7) ? 0 : this.y_value++;5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   U   c      3        = (this.y_value == 7) ? 0 : this.y_value++;5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   U   c      1        (this.y_value == 7) ? 0 : this.y_value++;5�_�   �   �           �   T   "    ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   V   c      3        if(this.y_value == 7) ? 0 : this.y_value++;5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   T   V   e                  �   T   V   d    5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   U   W   f              �   U   W   e    5�_�   �   �           �   W       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   V   X   f                  : this.y_value++;5�_�   �   �           �   W       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   V   X   f                   this.y_value++;5�_�   �   �           �   T       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   S   U   f              if(this.y_value == 7)5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   U   W   g                  �   U   W   f    5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   U   W   h                  �   U   W   g    5�_�   �   �           �   V       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   U   W   h                  if5�_�   �   �           �   V       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   U   W   h                  if()5�_�   �   �           �   V       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   U   W   h                  if()5�_�   �   �           �   V   !    ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   U   W   h      !            if(this.x_value == 7)5�_�   �   �           �   V   %    ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   V   Y   i                      �   V   X   h    5�_�   �   �           �   W        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   V   X   j       5�_�   �   �           �   X       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�    �   X   Z   k                  �   X   Z   j    5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   R   T   k          function getratio();5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   R   T   k          function getratiopair();5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5    �   R   T   k          function updatepair();5�_�   �   �           �   ]       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5    �   ]   _   k    5�_�   �   �           �   ^        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5     �   ]   ^           5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5&     �   F   H   k      6        !(size_in inside{no_size_inf, 'd5, 'd6, 'd7});5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5(     �   F   H   k      5        (size_in inside{no_size_inf, 'd5, 'd6, 'd7});5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5,     �   F   H   k      ,        (size_in inside{dl, 'd5, 'd6, 'd7});5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5.     �   F   H   k              (size_in inside{5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z52     �   F   H   k              (size_in inside{};5�_�   �   �           �   G       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5;    �   F   H   k              size_in inside{};5�_�   �   �           �   >        ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5H     �   =   >           5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   J   L   j          logic [2:0] x_value;5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�     �   K   L              logic [2:0] y_value;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�   	 �   J   L   i          logic [5:0] x_value;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            6   %       8          V   %    Z5�   
 �   J   L   i          logic [5:0] ratio_pair;5�_�   �   �           �   Q        ����                                                                                                                                                                                                                                                                                                                            Q   	       [   	       V   	    Z5�     �   P   Q              function updateRatioPair();   "        if(this.y_value == 7)begin               this.y_value = 0;   &            if(this.x_value == 7)begin   !                this.x_value = 0;               end               this.x_value++;           end           else                this.y_value++;       endfunction5�_�   �   �           �   L        ����                                                                                                                                                                                                                                                                                                                            Q   	       Q   	       V   	    Z5�     �   K   L              function new();5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            P   	       P   	       V   	    Z5�     �   K   L                  this.x_value = 0;5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            O   	       O   	       V   	    Z5�     �   K   L                  this.y_value = 0;5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            N   	       N   	       V   	    Z5�     �   K   L              endfunction5�_�   �   �           �   K        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   K   O   Z    �   K   L   Z    5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   N   P   ^          �   N   P   ]    5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   N   O              5�_�   �   �           �   O        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5    �   N   O           5�_�   �   �           �   X       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5]     �   W   Y   \              interval inside{1};5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5a     �   Z   _   ]       �   Z   \   \    5�_�   �   �           �   [        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5p     �   [   a   `    �   [   \   `    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5�    �         e      class supply_rand;5�_�   �   �           �   a        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5R     �   a   e   e    �   a   b   e    5�_�   �   �           �   d       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5�     �   c   e   h      flavor machine_flavor_out;5�_�   �   �           �   d   +    ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5�    �   c   e   h      2flavor machine_flavor_out;// To Compare The Output5�_�   �   �           �   d   %    ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5�     �   d   h   i       �   d   f   h    5�_�   �   �           �   g        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5�     �   f   h   k       5�_�   �   �           �   k       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z53     �   j              
endprogram5�_�   �   �           �   g        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   f   g          task 5�_�   �   �           �   f        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   f   h   k       �   f   h   j    5�_�   �   �           �   f        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5	     �   e   g   k       5�_�   �   �           �   h        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   h   j   l          �   h   j   k    5�_�   �   �           �   g       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   g   i   m          �   g   i   l    5�_�   �   �           �   h   	    ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   g   i   m      	    reset5�_�   �   �           �   h   
    ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5     �   g   i   m          reset()5�_�   �   �           �   l        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z5/     �   l   �   m    �   l   m   m    5�_�   �   �           �   o        ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z53     �   n   o          *    $display("*************************");5�_�   �   �           �   p       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z54     �   o   p          *    $display("*************************");5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                            A           C           V        Z58     �   l   n   �      task reset();    begin5�_�   �   �           �   x        ����                                                                                                                                                                                                                                                                                                                            x          �          V       Z5M     �   w   x              if((inf.out_valid !== 0)   )        || (inf.flavor_out !== no_coffee)   ,        || (inf.window.espresso.led !== red)   2        || (inf.window.espresso.monitor !== 10'd0)   (        || (inf.window.milk.led !== red)   .        || (inf.window.milk.monitor !== 10'd0)   -        || (inf.window.chocolate.led !== red)   3        || (inf.window.chocolate.monitor !== 10'd0)   )        || (inf.window.froth.led !== red)   /        || (inf.window.froth.monitor !== 10'd0)       )5�_�   �   �           �   w        ����                                                                                                                                                                                                                                                                                                                            x          x          V       Z5N     �   w   y   x    5�_�   �   �           �   w       ����                                                                                                                                                                                                                                                                                                                            y          y          V       Z5g     �   w   �   y    �   w   x   y    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5k     �   �   �          *    $display("*************************");5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5l     �   �   �          *    $display("*************************");5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5s     �   �   �   �    �   �   �   �    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5u     �   �   �   �       �   �   �   �    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5�     �   �   �   �      task input_supply5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5�     �   �   �   �      task input_supply()5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5y     �   �     �    �   �   �   �    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                              V       Z5~    �   �   �        task input_supply();5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                              V       Z5$    �   �   �        task input_supply(full);5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                              V       Z5F    �   �   �        5task input_supply(full); //policy always fill to full5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                                              V       Z5L     �   �   �        4task input_supply(full);//policy always fill to full5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                              V       Z5M    �   �   �         �   �   �      5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                              V       Z5�     �  
             5�_�   �   �           �  
       ����                                                                                                                                                                                                                                                                                                                                              V       Z5�     �  
              �  
        5�_�   �   �           �  
       ����                                                                                                                                                                                                                                                                                                                                              V       Z5�    �  
              �  
        5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                              V       Z5�    �   �   �        task input_supply(full);   begin5�_�   �   �           �         ����                                                                                                                                                                                                                                                                                                                                              V       Z5
     �             �          5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                              V       Z5    �    �      �          5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �      �      3task press_buttom(select_flavor select_flavor_rand,   /                  select_size select_size_rand,5�_�   �   �           �     3    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �      �      Qtask press_buttom(select_flavor select_flavor_rand, select_size select_size_rand,   2                  select_ratio select_ratio_rand);5�_�   �   �           �     Q    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5    �      �      rtask press_buttom(select_flavor select_flavor_rand, select_size select_size_rand, select_ratio select_ratio_rand);   begin5�_�   �   �   �       �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �              repeat(1)@(negedge clk);5�_�   �   �           �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �              out_valid_check();5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �              window_check();5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �              flavor_out_check();5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �              out_valid_one_cycle();5�_�   �   �           �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �           5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �              // after press button5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �  �  �          #    machine_flavor_out = no_coffee;5�_�   �   �           �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          task out_valid_check(); begin5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5
     �  �  �              check_output_times = 0;5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5
     �  �  �          ?    while(inf.out_valid !== 1 && check_output_times < 30) begin5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          -	check_output_times = check_output_times + 1;5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          	repeat(1)@(negedge clk);5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �              end5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          &    if(check_output_times == 30) begin5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          E	$display("-----Your out_valid should be high in 30 cycles------\n");5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �                  fail;5�_�   �   �           �  �       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �              end5�_�   �   �           �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          end5�_�   �   �           �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          endtask5�_�   �   �           �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �          ,//-----------Checkt out_valid---------------5�_�   �      �       �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5    �  �  �           5�_�   �                h       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5"     �   h   j  �          �   h   j  �    5�_�                  i       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5&     �   h   j  �          for 5�_�                 i   	    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5&     �   h   j  �      
    for ()5�_�                 i       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z58     �   h   j  �          for5�_�                 i       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z58     �   h   j  �      	    for()5�_�                 i       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5:     �   h   j  �      	    for()5�_�                 i   5    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5L     �   h   j  �      5    for(index_i = 0 ; index_i <  ; index = index + 1)5�_�                 i   9    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5N     �   i   k  �              �   i   k  �    5�_�    	             i       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5O     �   i   k  �    5�_�    
          	   j        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5b     �   i   k  �       5�_�  	            
   i        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   h   j  �      :    for(index_i = 0 ; index_i <  ; index = index + 1)begin5�_�  
             i   ;    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�    �   h   j  �      ;    for(index_i = 0 ; index_i < 5 ; index = index + 1)begin5�_�                 i   D    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �   i   k  �              �   i   k  �    5�_�                 j       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �   i   k  �              for5�_�                 j       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �   i   k  �              for()5�_�                 j       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �   i   k  �              for()5�_�                 j   P    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5+     �   i   k  �      P        for(index_flavor = 0; index_flavor < 3 ; index_flavor = index_flavor +1)5�_�                 j   T    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5,     �   j   l  �                  �   j   l  �    5�_�                 j   
    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5-     �   j   l  �    5�_�                 m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5.     �   l   m                  5�_�                 m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z50    �   m   o  �    5�_�                 j       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5C     �   j   l  �                  �   j   l  �    5�_�                 k       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5D     �   j   l  �                  for5�_�                 k   0    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5T     �   j   l  �      1            for(index_size = 0 ; index_size < 4;)5�_�                 k   0    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5U     �   j   l  �      1            for(index_size = 0 ; index_size < 4;)5�_�                 k   L    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5g     �   j   l  �      L            for(index_size = 0 ; index_size < 4; index_size = index_size +1)5�_�                 k   P    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5h     �   k   m  �                      �   k   m  �    5�_�                 l       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5j     �   k   m  �                      endk5�_�                 k       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5j     �   k   m  �    5�_�                 n        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5k     �   m   n           5�_�                  m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5m     �   l   n  �                      end5�_�    !              m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5n     �   l   n  �                 end5�_�     "          !   m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5n    �   l   n  �                 end5�_�  !  #          "   l        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   k   m  �       5�_�  "  $          #   l       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   k   m  �                      5�_�  #  %          $   l       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   k   m  �                      supply_input5�_�  $  &          %   l       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   k   m  �                      supply_input()5�_�  %  '          &   l       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   k   m  �                      supply_input()5�_�  &  (          '   l       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   k   m  �                      supply_input(1)5�_�  '  )          (   l   &    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   l   n  �    5�_�  (  *          )   l       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   l   n  �                      �   l   n  �    5�_�  )  +          *   m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   l   n  �                      press_buttom5�_�  *  ,          +   m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   l   n  �                      press_buttom()5�_�  +  -          ,   m       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   l   n  �                      press_buttom()5�_�  ,  .          -   m   D    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �   l   n  �      D                press_buttom(select_flavor_rand, select_size_rand,0)5�_�  -  /          .   m   C    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5    �   l   n  �      E                press_buttom(select_flavor_rand, select_size_rand,0);5�_�  .  0          /   m   R    ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5E     �   m   p  �    �   m   n  �    5�_�  /  1          0   n       ����                                                                                                                                                                                                                                                                                                                            n          o                 Z5I     �   m   p  �      9                        void'(interval_rand.randomize());   E                        repeat(interval_rand.interval)@(negedge clk);5�_�  0  2          1   l       ����                                                                                                                                                                                                                                                                                                                            n          o                 Z5K     �   l   n  �    5�_�  1  3          2  �        ����                                                                                                                                                                                                                                                                                                                            o          p                 Z5�     �  �  �  �    �  �  �  �    5�_�  2  4          3   n       ����                                                                                                                                                                                                                                                                                                                            o          p                 Z5�     �   n   p  �                      �   n   p  �    5�_�  3  5          4   o       ����                                                                                                                                                                                                                                                                                                                            p          q                 Z5�     �   o   q  �                      �   o   q  �    5�_�  4  6          5   n       ����                                                                                                                                                                                                                                                                                                                            q          r                 Z5�     �   n   p  �                      �   n   p  �    5�_�  5  7          6   o       ����                                                                                                                                                                                                                                                                                                                            r          s                 Z5�     �   n   p  �                      @5�_�  6  8          7   o   #    ����                                                                                                                                                                                                                                                                                                                            r          s                 Z5�     �   n   p  �      $                @(posedge out_valid)5�_�  7  9          8   o   $    ����                                                                                                                                                                                                                                                                                                                            r          s                 Z5�     �   n   p  �      $                @(posedge out_valid)5�_�  8  :          9   o   $    ����                                                                                                                                                                                                                                                                                                                            r          s                 Z5�     �   n   p  �      %                @(posedge out_valid);5�_�  9  ;          :   o   #    ����                                                                                                                                                                                                                                                                                                                            r          s                 Z5�    �   n   p  �      $                @(posedge out_valid)                   window_check;5�_�  :  <          ;   o       ����                                                                                                                                                                                                                                                                                                                            q          r                 Z5�     �   n   o          2                @(posedge out_valid) window_check;5�_�  ;  =          <   m        ����                                                                                                                                                                                                                                                                                                                            p          q                 Z5�     �   m   o  �    �   m   n  �    5�_�  <  >          =   m        ����                                                                                                                                                                                                                                                                                                                            q          r                 Z5�     �   l   m           5�_�  =  ?          >   m       ����                                                                                                                                                                                                                                                                                                                            p          q                 Z5�     �   m   p  �                      �   m   o  �    5�_�  >  @          ?   r        ����                                                                                                                                                                                                                                                                                                                            r          s          V       Z5�     �   q   r          1                void'(interval_rand.randomize());   =                repeat(interval_rand.interval)@(negedge clk);5�_�  ?  A          @   n        ����                                                                                                                                                                                                                                                                                                                            r          r          V       Z5�     �   n   q  �    �   n   o  �    5�_�  @  B          A   n        ����                                                                                                                                                                                                                                                                                                                            t          t          V       Z5�     �   m   n           5�_�  A  C          B   m       ����                                                                                                                                                                                                                                                                                                                            s          s          V       Z5�     �   m   o  �    5�_�  B  D          C   s        ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z5     �   s   v  �    �   s   t  �    5�_�  C  E          D   v        ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z5     �   u   v           5�_�  D  F          E   r       ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z5     �   r   t  �    �   r   s  �    5�_�  E  G          F   s   2    ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z5     �   r   t  �      2                @(posedge out_valid) window_check;5�_�  F  H          G  �       ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z5'     �  �  �  �    5�_�  G  I          H   s   3    ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z5+    �   r   t  �      3                @(posedge out_valid) window_check; 5�_�  H  J          I   t       ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z51     �   s   t                          5�_�  I  K          J   s       ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z52     �   s   u  �    5�_�  J  L          K   h       ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z55    �   h   j  �          �   h   j  �    5�_�  K  M          L  �        ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5X     �  �  +  �    �  �  �  �    5�_�  L  N          M   z       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5v     �   z   |  -          �   z   |  ,    5�_�  M  O          N  ,        ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  ,  f  -    �  ,  -  -    5�_�  N  P          O  /        ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          	repeat(10)@(negedge clk);5�_�  O  Q          P  /        ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /           5�_�  P  R          Q  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO");5�_�  Q  S          R  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOoooooo888888OOOOOOOOOOOOOOOOOOOOOOO");5�_�  R  T          S  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOO88OOoc:.                   cOOOOOOOOOOOOOOOOOOOOOOOOOOOOO");5�_�  S  U          T  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOOOOOOOOOOOOO8O.                             oOOOOOOOOOOOOOOOOOOOOOOOOOOOO");5�_�  T  V          U  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOOOOOOOOO8O.                                     oOOOOOOOOOOOOOOOOOOOOOOOO");5�_�  U  W          V  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOOOOOOOO:                                            O8OOOOOOOOOOOOOOOOOOO");5�_�  V  X          W  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOOOO8c                                                 O8OOOOOOOOOOOOOOOOO");5�_�  W  Y          X  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOOOO8.                                                     O8OOOOOOOOOOOOOOO");5�_�  X  Z          Y  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOO8.                                                         8OOOOOOOOOOOOOO");5�_�  Y  [          Z  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOOOOc                                                            oOOOOOOOOOOOOO");5�_�  Z  \          [  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOOO8c                                                              C8OOOOOOOOOOO");5�_�  [  ]          \  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOO8                                                                 .OOOOOOOOOOO");5�_�  \  ^          ]  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOOOO.                                                                  c8OOOOOOOOO");5�_�  ]  _          ^  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOO8                                                                      8OOOOOOOO");5�_�  ^  `          _  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOOOO:                      C.            :.            O@                  o8OOOOOOO");5�_�  _  a          `  /       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  .  /          e	$display("OOOOO8.                      O@@C          o@@8:        C@@@@C                 oOOOOOOO");5�_�  `  b          a  I       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  H  I          e	$display("OOOOOOOOOOOOOOO.   c@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:      COOOOOOOOOOOOO");5�_�  a  c          b  I       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  H  I          e	$display("OOOOOOOOOOOOOOOOOo    8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@O    O@8c  C8OOOOOOOOOOO");5�_�  b  d          c  I       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  H  I          e	$display("OOOOOOOOOOOOOOOOOOC.      O@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@8C     c@C  @8:   OOOOOOOOOOO");5�_�  c  e          d  I       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  H  I          e	$display("OOOOOOOOOOOOOOOOO8  .8         .oO@@@@@@@@@@@@@@@@@@8O:      c888888o  C8O  :8OOOOOOOOO");5�_�  d  f          e  I       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  H  I          e	$display("OOOOOOOOOOOOOOOO8c  88 .  ....                          oO888888888888  88c   8OOOOOOOO");5�_�  e  g          f  I       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  H  I          e	$display("OOOOOOOOOOOOOOOO.   @:.8.   ....  C@@8OOoocccoooO888888888888888888888O  C@C  8OOOOOOOO");5�_�  f  h          g  I        ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  H  I           5�_�  g  i          h  H       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5     �  G  H          e	$display("OOOOOOOOOOOOC    o@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@o   .COOOOOOOOOOOOO");   	$display("fail");5�_�  h  j          i  J       ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5   ! �  J  L  K    5�_�  i  k          j   e        ����                                                                                                                                                                                                                                                                                                                            p          q          V       Z5�     �   e   y  L    �   e   f  L    5�_�  j  l          k   i       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5�     �   h   j  _      int iter_i;5�_�  k  m          l   j       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5�     �   i   k  _      int iter_j;5�_�  l              m   k   
    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z5�   " �   j   l  _      int iter_k;5�_�  
               i       ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5�     �   h   j  �      7    for(ite = 0 ; index_i < 5 ; index = index + 1)begin5�_�   �           �   �  �        ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �  �  �        5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                           �         �          V       Z5     �            5�_�   �           �   �   �        ����                                                                                                                                                                                                                                                                                                                                              V       Z5I     �   �   �        5�_�   $           &   %   '       ����                                                                                                                                                                                                                                                                                                                            !   '       $                 Z5     �   '   (   +    �   &   ,          0            espresso_addnespresso_addnum;um > 0;   %        }                milk_addnum;   )endclass                 chocolate_addnum   )                         froth_addnum;      
endprogram5��