Vim�UnDo� � 2��طe'?X�#:b�j�
 ����sKq^��   �           2   v  ^  ^  �  ^  ]    Z4��    _�       w           v   <        ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2�V     �   ;   =   @      mEach combination should be pressed at least 5 times.((latte, cappuccino, mocha, user_define) x (s, m, l, xl))5�_�   v   x           w   =       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2�Y     �   =   ?   A          //�   =   ?   @    5�_�   w   y           x   >       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   =   ?   A      ,    cross cov_flavor_btn, cov_required_size;5�_�   x   z           y   =        ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   <   >   A          //cross coverage5�_�   y   {           z   >       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   >   @   B          �   >   @   A    5�_�   z   |           {   >       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   >   @   B    5�_�   {   }           |   >       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2�8     �   >   @   D          �   >   @   C    5�_�   |   ~           }   ?       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   ?   A   E          �   ?   A   D    5�_�   }              ~   >       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��    �   >   @   E    5�_�   ~   �              B        ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2�m     �   A   B           5�_�      �           �   C        ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2�p     �   C   E   F       �   C   E   E    5�_�   �   �           �   D       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2�{     �   C   E   F      covergroup cov_led @5�_�   �   �           �   D   !    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2�     �   C   E   F      !covergroup cov_led @(posedge clk)5�_�   �   �           �   D   !    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   F   G          �   D   F   F    5�_�   �   �           �   D       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   C   F   H      "covergroup cov_led @(posedge clk);    �   D   F   H          �   D   F   G    5�_�   �   �           �   E   /    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   F   H      ///Every ingredients’ led should be available 5�_�   �   �           �   E   5    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   F   H      6//Every ingredients’ led should be available (green)5�_�   �   �           �   E   L    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   H   H      L//Every ingredients’ led should be available (green) at least 1000 times. 5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   F   H   J      //inf.out_valid is high)5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   E   G   J      //(sample the value when   //inf.out_valid is high)5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   E   G   I      1//(sample the value when //inf.out_valid is high)5�_�   �   �           �   E       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   F   I      K//Every ingredients’ led should be available (green) at least 1000 times.   ///(sample the value when inf.out_valid is high)5�_�   �   �           �   E   L    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   F   H      |//Every ingredients’ led should be available (green) at least 1000 times.  //(sample the value when inf.out_valid is high)5�_�   �   �           �   E   L    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   F   H      {//Every ingredients’ led should be available (green) at least 1000 times. //(sample the value when inf.out_valid is high)5�_�   �   �           �   E   L    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   D   F   H      x//Every ingredients’ led should be available (green) at least 1000 times. sample the value when inf.out_valid is high)5�_�   �   �           �   E   L    ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   E   N   I      //�   E   G   H    5�_�   �   �           �   M       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   M   O   P    5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   E   G   Q          window.espresso.led green5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   E   G   Q          .espresso.led green5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   E   G   Q          espresso.led green5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   F   G              window.espresso.monitor 425�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   F   H   P          window.milk.led green5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          <           <   +          +    Z2��     �   F   H   P          .milk.led green5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          H          L   
          
    Z2��     �   G   M   P          window.milk.monitor 76       window.chocolate.led green        window.chocolate.monitor 110       window.froth.led green       windowsfroth.monito5�_�   �   �           �   L       ����                                                                                                                7                                                                                                                                                                                                          H          L   
          
    Z2��     �   K   L              froth.monito5�_�   �   �           �   J        ����                                                                                                                7                                                                                                                                                                                                          H          L   
          
    Z2��     �   I   J              chocolate.monitor 1105�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          H          K   
          
    Z2��     �   G   H              milk.monitor 765�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2��     �   F   H   M          milk.led green5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2��     �   G   I   M          chocolate.led green5�_�   �   �           �   I   	    ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2��     �   H   J   M          froth.led green5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�     �   E   G   M          espresso_led green5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�     �   E   G   M          espresso_ledgreen5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�
     �   F   H   M          milk_led green5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�     �   G   I   M          chocolate_led green5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�     �   G   I   M          chocolate_led g5�_�   �   �           �   I       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�     �   H   J   M          froth_led green5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�     �   E   G   M          espresso_led5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          H          J   
          
    Z2�     �   E   G   M          espresso_led 5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          F          I                 Z2�     �   E   G   M          espresso_led  5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          F          H                 Z2�      �   F   I   M          milk_led        chocolate_led �   E   G   M          espresso_led  5�_�   �   �           �   I       ����                                                                                                                7                                                                                                                                                                                                          F          H                 Z2�#     �   H   J   M          froth_led5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          F          H                 Z2�*     �   E   G   M          espresso_led  :5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          F          H                 Z2�8     �   F   H   M          milk_led      :5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          F          H                 Z2�;     �   F   H   M          milk_led      :P5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          F          H                 Z2�<     �   F   H   M          milk_led      :P{}5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          H          I                 Z2�l     �   G   I   M          chocolate_led :5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          H          I                 Z2�m     �   H   J   M          froth_led     :�   G   I   M          chocolate_led : 5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          H          I                 Z2�u     �   F   H   M          milk_led      :{}5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          H          I                 Z2�y     �   F   H   M          milk_led      : {}�   G   H   M    5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   F   K   M      &    milk_led      : {inf.window. .led}   &    chocolate_led : {inf.window. .led}   &    froth_led     : {inf.window. .led}    �   G   H   M    5�_�   �   �           �   G   (    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   F   H   M      3    milk_led      : {inf.window.milk_led      .led}5�_�   �   �           �   H   -    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   G   I   M      3    chocolate_led : {inf.window.chocolate_led .led}5�_�   �   �           �   I   )    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   H   J   M      3    froth_led     : {inf.window.froth_led     .led}5�_�   �   �           �   F   ,    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   E   G   M      ,    espresso_led  :{inf.window.espresso.led}5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   E   G   M      -    espresso_led  :{inf.window.espresso.led};5�_�   �   �           �   G   -    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   F   H   M      -    milk_led      : {inf.window.milk_led.led}5�_�   �   �           �   H   2    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   G   I   M      2    chocolate_led : {inf.window.chocolate_led.led}5�_�   �   �           �   H   .    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   G   I   M      3    chocolate_led : {inf.window.chocolate_led.led};5�_�   �   �           �   H   -    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   G   I   M      0    chocolate_led : {inf.window.chocolate_led.};5�_�   �   �           �   H   )    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   G   I   M      /    chocolate_led : {inf.window.chocolate_led};5�_�   �   �           �   G   $    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   F   H   M      .    milk_led      : {inf.window.milk_led.led};5�_�   �   �           �   I   %    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   H   J   M      .    froth_led     : {inf.window.froth_led.led}5�_�   �   �           �   I   *    ����                                                                                                                7                                                                                                                                                                                                          G          I                 Z2��     �   H   J   M      *    froth_led     : {inf.window.froth.led}5�_�   �   �           �   K       ����                                                                                                                7                                                                                                                                                                                                          @          @          V   *    Z2��     �   K   M   M    �   K   L   M    5�_�   �   �   �       �   F       ����                                                                                                                7                                                                                                                                                                                                          6          9                 Z2��     �   E   K   N      .    espresso_led  : {inf.window.espresso.led};   *    milk_led      : {inf.window.milk.led};   /    chocolate_led : {inf.window.chocolate.led};   +    froth_led     : {inf.window.froth.led};    �   F   G   N    5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          F          I                 Z2��     �   F   J   N      .    milk_led      : {binsinf.window.milk.led};   3    chocolate_led : {binsinf.window.chocolate.led};   /    froth_led     : {binsinf.window.froth.led};�   E   G   N      2    espresso_led  : {binsinf.window.espresso.led};5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          F          I                 Z2��     �   E   H   N      3    espresso_led  : {bins inf.window.espresso.led};5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          F          J                 Z2��     �   G   I   O      /    milk_led      : {bins inf.window.milk.led};5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          F          J                 Z2��     �   G   J   O      /    milk_led      : {bins inf.window.milk.led};5�_�   �   �           �   J       ����                                                                                                                7                                                                                                                                                                                                          F          K                 Z2��     �   I   L   P      4    chocolate_led : {bins inf.window.chocolate.led};5�_�   �   �           �   L       ����                                                                                                                7                                                                                                                                                                                                          F          L                 Z2��     �   K   N   Q      0    froth_led     : {bins inf.window.froth.led};5�_�   �   �           �   G   %    ����                                                                                                                7                                                                                                                                                                                                          F          L                 Z2�     �   F   H   R      &        bins inf.window.espresso.led};5�_�   �   �           �   G   (    ����                                                                                                                7                                                                                                                                                                                                          F          L                 Z2�     �   F   H   R      )        bins inf.window.espresso.led} = ;5�_�   �   �           �   G   )    ����                                                                                                                7                                                                                                                                                                                                          F          L                 Z2�     �   F   H   R      +        bins inf.window.espresso.led} = {};5�_�   �   �           �   G   )    ����                                                                                                                7                                                                                                                                                                                                          F          L                 Z2�     �   F   H   R      +        bins inf.window.espresso.led} = {};5�_�   �   �           �   G   0    ����                                                                                                                7                                                                                                                                                                                                          F          L                 Z2�     �   F   J   R      0        bins inf.window.espresso.led} = {green};5�_�   �   �           �   I        ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�     �   H   J   T      }5�_�   �   �           �   H        ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�     �   G   I   T       5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�"     �   G   I   T              bins ignore_bins5�_�   �   �           �   H       ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�(     �   G   I   T              ignore_bins5�_�   �   �           �   G   $    ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�2     �   F   H   T      0        bins inf.window.espresso.led} = {green};5�_�   �   �           �   H   "    ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�4     �   G   I   T      "        ignore_bins espresso_red =5�_�   �   �           �   H   #    ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�5     �   G   I   T      #        ignore_bins espresso_red = 5�_�   �   �           �   H   (    ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�7     �   G   I   T      (        ignore_bins espresso_red = {red}5�_�   �   �           �   K   !    ����                                                                                                                7                                                                                                                                                                                                          F          N                 Z2�;     �   K   M   T    �   K   L   T    5�_�   �   �           �   N       ����                                                                                                                7                                                                                                                                                                                                          F          O                 Z2�<     �   N   P   U    �   N   O   U    5�_�   �   �           �   Q       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�=     �   Q   S   V    �   Q   R   V    5�_�   �   �           �   Q   !    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�@     �   P   R   W      #        bins inf.window.froth.led};5�_�   �   �           �   Q   !    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�A     �   P   R   W      "        bins inf.window.froth.led;5�_�   �   �           �   Q   $    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�B     �   P   R   W      %        bins inf.window.froth.led = ;5�_�   �   �           �   Q   *    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�E     �   P   R   W      ,        bins inf.window.froth.led = {green};5�_�   �   �           �   N   %    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�G     �   M   O   W      '        bins inf.window.chocolate.led};5�_�   �   �           �   N   &    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�G     �   M   O   W      &        bins inf.window.chocolate.led;5�_�   �   �           �   N   (    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�L     �   M   O   W      )        bins inf.window.chocolate.led = ;5�_�   �   �           �   N   )    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�L     �   M   O   W      +        bins inf.window.chocolate.led = {};5�_�   �   �           �   N   )    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�M     �   M   O   W      +        bins inf.window.chocolate.led = {};5�_�   �   �           �   K        ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�P     �   J   L   W      "        bins inf.window.milk.led};5�_�   �   �           �   K   #    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�Q     �   J   L   W      %        bins inf.window.milk.led = };5�_�   �   �           �   K   )    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�S     �   J   L   W      ,        bins inf.window.milk.led = {green}};5�_�   �   �           �   K   *    ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�T     �   J   L   W      ,        bins inf.window.milk.led = {green}};5�_�   �   �           �   L       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�X     �   K   M   W      )        ignore_bins espresso_red = {red};5�_�   �   �           �   L       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�Z     �   K   M   W      "        ignore_bins o_red = {red};5�_�   �   �           �   O       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�f     �   N   P   W      )        ignore_bins espresso_red = {red};5�_�   �   �           �   O       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�f     �   N   P   W      !        ignore_bins _red = {red};5�_�   �   �           �   O       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�g     �   N   P   W      !        ignore_bins _red = {red};5�_�   �   �           �   R       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�k     �   Q   S   W      )        ignore_bins espresso_red = {red};5�_�   �   �           �   R       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�k     �   Q   S   W      !        ignore_bins _red = {red};5�_�   �   �           �   R       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�m     �   Q   S   W      !        ignore_bins _red = {red};5�_�   �   �           �   R       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�p     �   R   T   X              �   R   T   W    5�_�   �   �   �       �   O       ����                                                                                                                7                                                                                                                                                                                                          F          P                 Z2�u     �   O   Q   Y              �   O   Q   X    5�_�   �   �           �   L       ����                                                                                                                7                                                                                                                                                                                                          F          Q                 Z2�w     �   L   N   Z              �   L   N   Y    5�_�   �   �           �   X       ����                                                                                                                7                                                                                                                                                                                                          F          R                 Z2��     �   X   Z   [          �   X   Z   Z    5�_�   �   �           �   V        ����                                                                                                                7                                                                                                                                                                                                          F          R                 Z2��     �   U   V           5�_�   �   �           �   X       ����                                                                                                                7                                                                                                                                                                                                          F          R                 Z2��     �   X   [   [       �   X   Z   Z    5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   F   H   \      /        bins inf.window.espresso.led = {green};5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   E   G   \          espresso_led  : {5�_�   �   �           �   F       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   E   H   \           espresso_led  :coverpoint  {           bins  = {green};�   F   G   \    5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   F   H   \              bins  = {green};5�_�   �   �           �   G       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   F   H   \      '        bins  espresso_green = {green};5�_�   �   �           �   J       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   I   K   \          milk_led      : {5�_�   �   �           �   K        ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   J   L   \      +        bins inf.window.milk.led = {green};5�_�   �   �           �   K        ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   J   L   \      +        bins inf.window.milk.led = {green};5�_�   �   �           �   K   !    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   J   L   \      -        bins inf.window.milk.led{} = {green};5�_�   �              �   K   "    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   J   M   \      -        bins inf.window.milk.led{} = {green};5�_�   �     �          J   
    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   I   K   ]          milk_led      :    !        bins inf.window.milk.led{5�_�                  J       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   I   K   \      -    milk_led      : bins inf.window.milk.led{5�_�                 J       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   I   K   \      (    milk_led      : inf.window.milk.led{5�_�                 K       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�     �   J   L   \                  = {green};5�_�                 N       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�$     �   M   O   \          chocolate_led : {5�_�                 N       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�$     �   M   O   \          chocolate_led :    0        bins inf.window.chocolate.led = {green};5�_�                 N       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�&     �   M   O   [      <    chocolate_led : bins inf.window.chocolate.led = {green};5�_�                 N       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�'     �   M   O   [      7    chocolate_led : inf.window.chocolate.led = {green};5�_�    	             N   6    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�,     �   M   O   [      A    chocolate_led :coverpoint inf.window.chocolate.led = {green};5�_�    
          	   N   6    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�,     �   M   O   [      A    chocolate_led :coverpoint inf.window.chocolate.led = {green};5�_�  	            
   N   7    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�-     �   M   O   [      C    chocolate_led :coverpoint inf.window.chocolate.led{} = {green};5�_�  
               N   8    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�-     �   M   O   [      C    chocolate_led :coverpoint inf.window.chocolate.led{} = {green};5�_�                 N   6    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�/     �   M   O   [      B    chocolate_led :coverpoint inf.window.chocolate.led{ = {green};5�_�                 N   8    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�0     �   M   P   [      C    chocolate_led :coverpoint inf.window.chocolate.led { = {green};5�_�                 R       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�?     �   Q   S   \          froth_led     : {5�_�                 R       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�A     �   Q   S   \          froth_led     :coverpoint {5�_�                 R       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�B     �   Q   S   \          froth_led     :coverpoint{5�_�                 R       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�C     �   Q   S   \          froth_led     :coverpoint   ,        bins inf.window.froth.led = {green};5�_�                 R       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�D     �   Q   S   [      B    froth_led     :coverpoint bins inf.window.froth.led = {green};5�_�                 R       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�E     �   Q   S   [      A    froth_led     :coverpointbins inf.window.froth.led = {green};5�_�                 R       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�I     �   Q   S   [      <    froth_led     :coverpointinf.window.froth.led = {green};5�_�                 R   2    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�M     �   Q   S   [      =    froth_led     :coverpoint inf.window.froth.led = {green};5�_�                 R   3    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�N     �   Q   S   [      >    froth_led     :coverpoint inf.window.froth.led  = {green};5�_�                 R   4    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�O     �   Q   S   [      @    froth_led     :coverpoint inf.window.froth.led {} = {green};5�_�                 R   5    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2�O    �   Q   T   [      @    froth_led     :coverpoint inf.window.froth.led {} = {green};5�_�                 D       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   C   E   \      "covergroup cov_led @(posedge clk);5�_�                 E       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   D   F   \      y//Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)5�_�                 E       ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   D   F   \      �    option.comment = Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)5�_�                 E   �    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   D   F   \      �    option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)5�_�                 ,        ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   +   ,          //  For Eazy to read5�_�                 +        ����                                                                                                                6                                                                                                                                                                                                          F          F   #          #    Z2��     �   *   ,   [      O//Every case of flavor_btn except no_coffee should be pressed at least 5 times.5�_�                  3        ����                                                                                                                6                                                                                                                                                                                                          F          F   #          #    Z2��     �   2   3          U//Every case of required_size expcept no_size_inf should be pressed at least 5 times.5�_�    !              +       ����                                                                                                                5                                                                                                                                                                                                          E          E   #          #    Z2��     �   +   -   Z    �   +   ,   Z    5�_�     "          !   ;        ����                                                                                                                6                                                                                                                                                                                                          F          F   #          #    Z2�      �   :   ;          o//Each combination should be pressed at least 5 times.((latte, cappuccino, mocha, user_define) x (s, m, l, xl))5�_�  !  #          "   ,        ����                                                                                                                6                                                                                                                                                                                                          E          E   #          #    Z2�     �   ,   .   Z    �   ,   -   Z    5�_�  "  $          #   <        ����                                                                                                                7                                                                                                                                                                                                          F          F   #          #    Z2�     �   ;   <          //cross coverage5�_�  #  %          $   -       ����                                                                                                                7                                                                                                                                                                                                          E          E   #          #    Z2�     �   -   /   Z    �   -   .   Z    5�_�  $  &          %   ,        ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   +   /   [      U//Every case of required_size expcept no_size_inf should be pressed at least 5 times.   o//Each combination should be pressed at least 5 times.((latte, cappuccino, mocha, user_define) x (s, m, l, xl))   //cross coverage5�_�  %  '          &   .       ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�
     �   -   /   [      cross coverage5�_�  &  (          '   .       ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   -   /   [      cross coverage5�_�  '  )          (   +       ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   *   ,   [      MEvery case of flavor_btn except no_coffee should be pressed at least 5 times.5�_�  (  *          )   +        ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   *   ,   [      MEvery case of flavor_btn except no_coffee should be pressed at least 5 times.5�_�  )  +          *   +        ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   *   ,   [      N"Every case of flavor_btn except no_coffee should be pressed at least 5 times.5�_�  *  ,          +   +       ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   *   ,   [      _option.comment = "Every case of flavor_btn except no_coffee should be pressed at least 5 times.5�_�  +  -          ,   .       ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   -   /   [      cross coverage"5�_�  ,  .          -   +   ^    ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�     �   *   ,   [      ^option.comment ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.5�_�  -  /          .   ,   S    ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�"     �   +   -   [      SEvery case of required_size expcept no_size_inf should be pressed at least 5 times.5�_�  .  0          /   -   m    ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�$     �   ,   .   [      mEach combination should be pressed at least 5 times.((latte, cappuccino, mocha, user_define) x (s, m, l, xl))5�_�  /  1          0   .       ����                                                                                                                8                                                                                                                                                                                                          ,           .                 Z2�'     �   .   0   [    5�_�  0  2          1   X        ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�2     �   X   [   ]       �   X   Z   \    5�_�  1  3          2   .        ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�_     �   .   0   _       �   .   0   ^    5�_�  2  4          3   /        ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2�e     �   .   /          option.goal = 5;5�_�  3  5          4   ?        ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�i     �   ?   A   ^    �   ?   @   ^    5�_�  4  6          5   @       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�i     �   ?   A   _      option.goal = 5;5�_�  5  7          6   @        ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�j     �   ?   A   _      option.goal = 5;5�_�  6  8          7   @       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�o    �   ?   @              option.goal = 5;5�_�  7  9          8   Y        ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   X   [   ^       5�_�  8  :          9   Z       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   Y   [   _      covergroup cg_ratio_tran @5�_�  9  ;          :   Z   '    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   Y   [   _      'covergroup cg_ratio_tran @(posedge clk)5�_�  :  <          ;   Z   '    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   Z   ]   `          �   Z   \   _    5�_�  ;  =          <   Z       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   Z   \   b          �   Z   \   a    5�_�  <  >          =   [       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   Z   \   b          option.comment = 5�_�  =  ?          >   S       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   R   T   b      +        bins        froth_green  = {green};5�_�  >  @          ?   E   �    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   D   F   b      �    option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)"5�_�  ?  A          @   [       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   Z   ]   b          option.comment = "";5�_�  @  B          A   \   7    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   \   ^   d       �   \   ^   c    5�_�  A  C          B   ]       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   \   `   d          ratio_train : 5�_�  B  D          C   _       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ^   `   f          }5�_�  C  E          D   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�      �   ]   _   f          5�_�  D  F          E   ]       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�/     �   \   ^   f          ratio_train : {5�_�  E  H          F   ]       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�0     �   \   ^   f          ratio_tran : {5�_�  F  I  G      H   0       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�H     �   /   1   f      /    cov_flavor_btn: coverpoint inf.flavor_btn{ 5�_�  H  J          I   0       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�J     �   /   1   f      +    flavor_btn: coverpoint inf.flavor_btn{ 5�_�  I  K          J   7       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�P     �   6   8   f      4    cov_required_size: coverpoint inf.required_size{5�_�  J  L          K   7       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�R     �   6   8   f      0    required_size: coverpoint inf.required_size{5�_�  K  M          L   >       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�W     �   =   ?   f      ?    cross_cov_btn_size:cross cov_flavor_btn, cov_required_size;5�_�  L  N          M   F       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�d     �   E   G   f      7    espresso_led  :coverpoint inf.window.espresso.led {5�_�  M  O          N   J       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�h     �   I   K   f      3    milk_led      :coverpoint  inf.window.milk.led{5�_�  N  P          O   N       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�l     �   M   O   f      8    chocolate_led :coverpoint inf.window.chocolate.led {5�_�  O  Q          P   R       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�q     �   Q   S   f      4    froth_led     :coverpoint inf.window.froth.led {5�_�  P  R          Q   R       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�t    �   Q   S   f      7    froth_led_cpt    :coverpoint inf.window.froth.led {5�_�  Q  S          R   ]       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�z     �   \   ^   f          ratio_transition : {5�_�  R  T          S   ]       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              �   ]   _   f    5�_�  S  U          T   ]       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   \   ^   g          ratio_transition_cpt : {5�_�  T  V          U   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins 5�_�  U  W          V   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr5�_�  V  X          W   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[]5�_�  W  Y          X   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = 5�_�  X  Z          Y   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {}5�_�  Y  [          Z   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {[]}5�_�  Z  \          [   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {[]}5�_�  [  ]          \   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {[]}5�_�  \  ^          ]   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {[0:7]}5�_�  ]  _          ^   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {[0:7],}5�_�  ^  `          _   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {[0:7],[]}5�_�  _  a          `   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g              bins tr[] = {[0:7],[]}5�_�  `  b          a   ^       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g      !        bins tr[] = {[0:7],[0:7]}5�_�  a  c          b   ^   $    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ]   _   g      $        bins tr[] = {[0:7] => [0:7]}5�_�  b  d          c   _       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2��     �   ^   `   g              5�_�  c  e          d   _   #    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�     �   ^   `   g      #        bins other_trans = default;5�_�  d  f          e   <   .    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�;     �   ;   =   g      L        ignore_bins size_bad    = default; // each coverpoint is independent5�_�  e  g          f   <   .    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�<     �   ;   =   g      G        ignore_bins size_bad    = default; // coverpoint is independent5�_�  f  h          g   <   .    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�=     �   ;   =   g      <        ignore_bins size_bad    = default; // is independent5�_�  g  i          h   <   +    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�>     �   ;   =   g      .        ignore_bins size_bad    = default; // 5�_�  h  j          i   <   +    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�>     �   ;   =   g      -        ignore_bins size_bad    = default; / 5�_�  i  k          j   <   )    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�O     �   ;   =   g      ,        ignore_bins size_bad    = default;  5�_�  j  l          k   <   "    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�Q     �   ;   =   g      %        ignore_bins size_bad    = ;  5�_�  k  m          l   <   .    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�X     �   ;   =   g      2        ignore_bins size_bad    = {no_size_inf};  5�_�  l  n          m   5   !    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�]     �   4   6   g      *        ignore_bins btn_bad     = default;5�_�  m  o          n   5   "    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�^     �   4   6   g      #        ignore_bins btn_bad     = ;5�_�  n  p          o   5   ,    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�a     �   4   6   g      .        ignore_bins btn_bad     = {no_coffee};5�_�  o  q          p   5   +    ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�a     �   5   7   h              �   5   7   g    5�_�  p  r          q   =       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2�k     �   =   ?   h    �   =   >   h    5�_�  q  s          r   =       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2�r     �   <   >   i      2        ignore_bins size_bad    = {no_size_inf};  5�_�  r  t          s   =       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2�u     �   <   >   i      &        ignore_bins = {no_size_inf};  5�_�  s  u          t   =       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2�y     �   <   >   i      1        ignore_bins no_size_bin= {no_size_inf};  5�_�  t  v          u   >       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2�|     �   =   ?   i              illegal_bins = default;5�_�  u  w          v   >       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2�~     �   =   ?   i               illegal_bins  = default;5�_�  v  x          w   6       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2��     �   5   7   i              illegal_bins = default;5�_�  w  y          x   5       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2��     �   4   6   i      .        ignore_bins btn_bad     = {no_coffee};5�_�  x  z          y   5       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2��     �   4   6   i      (        ignore_bins d     = {no_coffee};5�_�  y  {          z   5   $    ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2��     �   4   6   i      5        ignore_bins  no_coffee_bin     = {no_coffee};5�_�  z  |          {   a       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2��     �   `   b   i      >        bins other_trans = default;// should get error message5�_�  {  }          |   ^       ����                                                                                                                :                                                                                                                                                                                                          ,           .                 Z2��     �   ^   `   j       �   ^   `   i    5�_�  |  ~          }   X        ����                                                                                                                :                                                                                                                                                                                                          X          Y          V       Z2��     �   W   X              option.at_least = 1000;       option.per_instance = 1;5�_�  }            ~   G        ����                                                                                                                :                                                                                                                                                                                                          X          X          V       Z2��     �   G   J   h    �   G   H   h    5�_�  ~  �             I       ����                                                                                                                :                                                                                                                                                                                                          Z          Z          V       Z2��     �   I   K   j    5�_�    �          �   G       ����                                                                                                                :                                                                                                                                                                                                          G          I                 Z2��     �   F   H   k      �    option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   H       ����                                                                                                                :                                                                                                                                                                                                          G          I                 Z2��     �   G   I   k          option.at_least = 1000;5�_�  �  �          �   I       ����                                                                                                                :                                                                                                                                                                                                          G          I                 Z2��     �   H   J   k          option.per_instance = 1;5�_�  �  �          �   B        ����                                                                                                                :                                                                                                                                                                                                          B          C          V       Z2��     �   A   B              option.at_least = 5;       option.per_instance = 1;5�_�  �  �          �   .        ����                                                                                                                :                                                                                                                                                                                                          B          B          V       Z2��     �   .   1   i    �   .   /   i    5�_�  �  �          �   +       ����                                                                                                                <                                                                                                                                                                                                          D          D          V       Z2��     �   *   ,   k      `option.comment ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   +        ����                                                                                                                <                                                                                                                                                                                                          D          D          V       Z2��     �   *   ,   k      `option.comment ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   g        ����                                                                                                                <                                                                                                                                                                                                          D          D          V       Z2�     �   g   i   l       �   g   i   k    5�_�  �  �          �   h       ����                                                                                                                <                                                                                                                                                                                                          D          D          V       Z2�     �   h   j   m       �   h   j   l    5�_�  �  �          �   i       ����                                                                                                                <                                                                                                                                                                                                          D          D          V       Z2�     �   i   k   n       �   i   k   m    5�_�  �  �          �   j        ����                                                                                                                <                                                                                                                                                                                                          D          D          V       Z2�"     �   i   j          cg_btn_required_size_crossdd5�_�  �  �          �   i        ����                                                                                                                <                                                                                                                                                                                                          D          D          V       Z2�#     �   i   k   n       �   i   k   m    5�_�  �  �          �   h        ����                                                                                                                <                                                                                                                                                                                                          h          j          V       Z2�*     �   g   h          cg_btn_required_size_cross   cg_led   cg_ratio_tran5�_�  �  �          �   i        ����                                                                                                                <                                                                                                                                                                                                          h          h          V       Z2�,     �   i   m   k    �   i   j   k    5�_�  �  �          �   i        ����                                                                                                                <                                                                                                                                                                                                          h          h          V       Z2�,     �   h   i          covergroup 5�_�  �  �          �   i        ����                                                                                                                <                                                                                                                                                                                                          h          h          V       Z2�<     �   h   i          cg_btn_required_size_cross5�_�  �  �          �   h        ����                                                                                                                <                                                                                                                                                                                                          h          h          V       Z2�=     �   h   j   m       �   h   j   l    5�_�  �  �          �   i       ����                                                                                                                <                                                                                                                                                                                                          h          h          V       Z2�Q     �   h   j   m      cg_btn_size_cross5�_�  �  �          �   i   .    ����                                                                                                                <                                                                                                                                                                                                          h          h          V       Z2�\     �   h   j   m      .cg_btn_size_cross cg_btn_size_cross_inst = new5�_�  �  �          �   i   /    ����                                                                                                                <                                                                                                                                                                                                          h          h          V       Z2�\     �   h   j   m      0cg_btn_size_cross cg_btn_size_cross_inst = new()5�_�  �  �          �   j       ����                                                                                                                <                                                                                                                                                                                                          j           k                 Z2�c     �   i   k   m      cg_led5�_�  �  �          �   j       ����                                                                                                                <                                                                                                                                                                                                          j           k                 Z2�f     �   i   m   m      cg_led              cg_ratio_tran    �   j   k   m    5�_�  �  �          �   j       ����                                                                                                                <                                                                                                                                                                                                          j          k                 Z2�h     �   j   l   m      cg_ratio_tran    cg_ratio_tran�   i   k   m      cg_led           cg_led5�_�  �  �          �   j       ����                                                                                                                <                                                                                                                                                                                                          j          k                 Z2�k     �   i   k   m      cg_led            cg_led5�_�  �  �          �   j       ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2�q     �   i   k   m      (cg_led            cg_led                5�_�  �  �          �   j   .    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2�t     �   i   k   m      7cg_led            cg_led                 = new         5�_�  �  �          �   j   /    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2�w     �   i   k   m      9cg_led            cg_led                 = new()         5�_�  �  �          �   j   0    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2�x     �   j   l   m      cg_ratio_tran     cg_ratio_tran�   i   k   m      9cg_led            cg_led                 = new()         5�_�  �  �          �   j       ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��     �   i   k   m      :cg_led            cg_led                 = new();         5�_�  �  �          �   j   )    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��     �   i   k   m      ?cg_led            cg_led_inst                 = new();         5�_�  �  �          �   k       ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��     �   j   l   m      1cg_ratio_tran     cg_ratio_tran          = new();5�_�  �  �          �   k   !    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��     �   j   l   m      6cg_ratio_tran     cg_ratio_tran_isnt          = new();5�_�  �  �          �   k   "    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��     �   j   l   m      6cg_ratio_tran     cg_ratio_tran_innt          = new();5�_�  �  �          �   k   "    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��     �   j   l   m      6cg_ratio_tran     cg_ratio_tran_inrt          = new();5�_�  �  �          �   k   "    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��     �   j   l   m      5cg_ratio_tran     cg_ratio_tran_int          = new();5�_�  �  �          �   k   )    ����                                                                                                                <                                                                                                                                                                                                          j   '       k             '    Z2��    �   j   l   m      6cg_ratio_tran     cg_ratio_tran_inst          = new();5�_�  �  �          �   ^        ����                                                                                                                <                                                                                                                                                                                                          ^   )       `          V   )    Z2��     �   ]   ^          |    option.comment = "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit   :    at least 50 times. (sample the value at posedge clk)";       option.at_least = 50;5�_�  �  �          �   `       ����                                                                                                                <                                                                                                                                                                                                          ^   )       ^          V   )    Z2��     �   `   d   j    �   `   a   j    5�_�  �  �          �   a       ����                                                                                                                <                                                                                                                                                                                                          a          c                 Z2��     �   a   d   m      :    at least 50 times. (sample the value at posedge clk)";       option.at_least = 50;�   `   b   m      |    option.comment = "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit5�_�  �  �          �   ]        ����                                                                                                                <                                                                                                                                                                                                          a          c                 Z2��     �   \   ]          (covergroup cg_ratio_tran @(posedge clk);5�_�  �  �          �   ]       ����                                                                                                                <                                                                                                                                                                                                          `          b                 Z2��     �   \   ^   l      &    ratio_transition_cpt : inf.ratio {5�_�  �  �          �   [        ����                                                                                                                <                                                                                                                                                                                                          `          b                 Z2��     �   Z   [          endgroup5�_�  �  �          �   [        ����                                                                                                                <                                                                                                                                                                                                          _          a                 Z2��     �   Z   [           5�_�  �  �          �   Z       ����                                                                                                                <                                                                                                                                                                                                          ^          `                 Z2��     �   Z   \   j    5�_�  �  �          �   H        ����                                                                                                                <                                                                                                                                                                                                          H          I          V       Z2��     �   G   H             option.at_least = 1000;      option.per_instance = 1;5�_�  �  �          �   K        ����                                                                                                                <                                                                                                                                                                                                          H          H          V       Z2��     �   K   N   i    �   K   L   i    5�_�  �  �          �   L       ����                                                                                                                <                                                                                                                                                                                                          L          M                 Z2��     �   L   N   k         option.per_instance = 1;�   K   M   k         option.at_least = 1000;5�_�  �  �          �   Q        ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2��     �   Q   T   k    �   Q   R   k    5�_�  �  �          �   W        ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2��     �   W   Z   m    �   W   X   m    5�_�  �  �          �   ]       ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2��     �   ]   `   o    �   ]   ^   o    5�_�  �  �          �   G       ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2��     �   F   G          �   option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   H        ����                                                                                                                <                                                                                                                                                                                                          K          L          V       Z2��     �   H   J   p    �   H   I   p    5�_�  �  �          �   O       ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2�      �   O   Q   q    �   O   P   q    5�_�  �  �          �   I       ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2�     �   H   J   r      �   option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   I       ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2�     �   H   J   r      �   option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   P       ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2�     �   O   Q   r      �   option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   V        ����                                                                                                                <                                                                                                                                                                                                          P          P          V       Z2�     �   V   X   r    �   V   W   r    5�_�  �  �          �   ]       ����                                                                                                                <                                                                                                                                                                                                          P          P          V       Z2�     �   ]   _   s    �   ]   ^   s    5�_�  �  �          �   a        ����                                                                                                                <                                                                                                                                                                                                          a          b          V       Z2�"     �   `   a                  option.at_least = 1000;            option.per_instance = 1;5�_�  �  �          �   ^       ����                                                                                                                <                                                                                                                                                                                                          a          a          V       Z2�$     �   ^   a   r    �   ^   _   r    5�_�  �  �          �   W       ����                                                                                                                <                                                                                                                                                                                                          c          c          V       Z2�&     �   W   Z   t    �   W   X   t    5�_�  �  �          �   \        ����                                                                                                                <                                                                                                                                                                                                          \          ]          V       Z2�(     �   [   \                  option.at_least = 1000;            option.per_instance = 1;5�_�  �  �          �   P       ����                                                                                                                <                                                                                                                                                                                                          \          \          V       Z2�,     �   P   S   t    �   P   Q   t    5�_�  �  �          �   U       ����                                                                                                                <                                                                                                                                                                                                          ^          ^          V       Z2�-     �   T   U                  option.at_least = 1000;5�_�  �  �          �   U       ����                                                                                                                <                                                                                                                                                                                                          ]          ]          V       Z2�.     �   T   U                   option.per_instance = 1;5�_�  �  �          �   L        ����                                                                                                                <                                                                                                                                                                                                          L          M          V       Z2�0     �   K   L                  option.at_least = 1000;            option.per_instance = 1;5�_�  �  �          �   H       ����                                                                                                                <                                                                                                                                                                                                          L          L          V       Z2�5     �   H   K   r    �   H   I   r    5�_�  �  �          �   J       ����                                                                                                                <                                                                                                                                                                                                          N          N          V       Z2�\     �   I   J                   option.per_instance = 1;5�_�  �  �          �   Q       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2�_     �   P   Q                   option.per_instance = 1;5�_�  �  �          �   I       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2�a     �   H   I                  option.at_least = 1000;5�_�  �  �          �   I       ����                                                                                                                <                                                                                                                                                                                                          L          L          V       Z2�d     �   I   K   q    �   I   J   q    5�_�  �  �          �   W       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2�f     �   V   W                   option.per_instance = 1;5�_�  �  �          �   ]       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2�h     �   \   ]                   option.per_instance = 1;5�_�  �  �          �   F        ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2�o     �   E   F          !covergroup cg_led @(posedge clk);5�_�  �  �          �   D        ����                                                                                                                <                                                                                                                                                                                                          L          L          V       Z2�q     �   C   D          endgroup5�_�  �  �          �   B       ����                                                                                                                <                                                                                                                                                                                                          K          K          V       Z2�y     �   A   C   n      ?    cross_cov_btn_size:cross cov_flavor_btn, cov_required_size;5�_�  �  �          �   B       ����                                                                                                                <                                                                                                                                                                                                          K          K          V       Z2�{     �   A   D   n      ?    cross_cov_btn_size:cross cov_flavor_btn, cov_required_size;5�_�  �  �          �   C       ����                                                                                                                <                                                                                                                                                                                                          L          L          V       Z2�~     �   C   E   p          �   C   E   o    5�_�  �  �          �   D       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2��     �   C   E   p      }a5�_�  �  �          �   D        ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2��     �   C   E   p      }5�_�  �  �          �   /       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2��     �   .   /              option.at_least = 5;5�_�  �  �          �   1       ����                                                                                                                ;                                                                                                                                                                                                          L          L          V       Z2��     �   1   3   o    �   1   2   o    5�_�  �  �          �   2       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2��     �   1   3   p          option.at_least = 5;5�_�  �  �          �   2       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2��     �   1   3   p          option.at_least = 5;5�_�  �  �          �   :       ����                                                                                                                <                                                                                                                                                                                                          M          M          V       Z2��     �   :   <   p    �   :   ;   p    5�_�  �  �          �   C       ����                                                                                                                =                                                                                                                                                                                                          N          N          V       Z2��     �   C   E   q    �   C   D   q    5�_�  �  �          �   +        ����                                                                                                                =                                                                                                                                                                                                          +          .          V       Z2��     �   *   +          d    option.comment ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n   UEvery case of required_size expcept no_size_inf should be pressed at least 5 times.\n   oEach combination should be pressed at least 5 times.((latte, cappuccino, mocha, user_define) x (s, m, l, xl))\n   cross coverage";5�_�  �  �          �   -       ����                                                                                                                9                                                                                                                                                                                                          +          +          V       Z2��     �   -   2   n    �   -   .   n    5�_�  �  �  �      �   .       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   -   /   r      d    option.comment ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   .       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   -   /   r      ^    .comment ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   .       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   -   /   r      ]    comment ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   .       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   -   /   r      U    ="Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   .       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   -   /   r      T    "Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   .       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   -   /   r      V    //"Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   1       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   0   2   r      cross coverage";5�_�  �  �          �   1       ����                                                                                                                =                                                                                                                                                                                                          +          +          V       Z2��     �   0   2   r      cross coverage"*5�_�  �  �          �   .        ����                                                                                                                =                                                                                                                                                                                                          .          1          V       Z2��     �   -   .          V    /*"Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n   UEvery case of required_size expcept no_size_inf should be pressed at least 5 times.\n   oEach combination should be pressed at least 5 times.((latte, cappuccino, mocha, user_define) x (s, m, l, xl))\n   cross coverage"*/5�_�  �  �          �   ,        ����                                                                                                                9                                                                                                                                                                                                          .          .          V       Z2��     �   ,   1   n    �   ,   -   n    5�_�  �  �          �   -        ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   ,   .   r      V    /*"Every case of flavor_btn except no_coffee should be pressed at least 5 times.\n5�_�  �  �          �   K       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   L   r      �        option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   K       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   L   r      �        .comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   K       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   L   r      �        comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   K       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   L   r      �        = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   K       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   L   r      �        "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   K   �    ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   L   r      �        /*"Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   K   �    ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   L   r      �        /*"Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";*/5�_�  �  �          �   K       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   J   K          �        /*"Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)"*/5�_�  �  �          �   I        ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   I   K   q    �   I   J   q    5�_�  �  �          �   J        ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   I   K   r      �        /*"Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)"*/5�_�  �  �          �   Q        ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2��     �   P   Q          �        option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   V       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2�     �   U   V          �        option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   [       ����                                                                                                                =                                                                                                                                                                                                          2          2          V       Z2�     �   Z   [          �        option.comment = "Every ingredients’ led should be available (green) at least 1000 times. (sample the value when inf.out_valid is high)";5�_�  �  �          �   c        ����                                                                                                                =                                                                                                                                                                                                          c          d          V       Z2�     �   b   c          �        option.comment = "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit   >        at least 50 times. (sample the value at posedge clk)";5�_�  �  �          �   _        ����                                                                                                                =                                                                                                                                                                                                          c          c          V       Z2�     �   _   b   m    �   _   `   m    5�_�  �  �          �   `        ����                                                                                                                =                                                                                                                                                                                                          e          e          V       Z2�
     �   _   a   o      �        option.comment = "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit5�_�  �  �          �   `        ����                                                                                                                =                                                                                                                                                                                                          e          e          V       Z2�     �   _   a   o      xoption.comment = "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit5�_�  �  �          �   `        ����                                                                                                                =                                                                                                                                                                                                          e          e          V       Z2�     �   _   a   o      r.comment = "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit5�_�  �  �          �   `        ����                                                                                                                =                                                                                                                                                                                                          e          e          V       Z2�     �   _   a   o      qcomment = "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit5�_�  �  �          �   `        ����                                                                                                                =                                                                                                                                                                                                          e          e          V       Z2�     �   _   a   o      i= "Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit5�_�  �  �          �   `        ����                                                                                                                =                                                                                                                                                                                                          e          e          V       Z2�     �   _   a   o      g"Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit5�_�  �  �          �   `       ����                                                                                                                =                                                                                                                                                                                                          e          e          V       Z2�     �   _   a   o      i//"Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit   >        at least 50 times. (sample the value at posedge clk)";5�_�  �  �          �   `       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�     �   _   a   n      �//"Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit at least 50 times. (sample the value at posedge clk)";5�_�  �  �          �   `   �    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�     �   _   a   n      �/*"Create the transitions bin for the inf.ratio signal from [0:7] to [0:7]. Each transition should be hit at least 50 times. (sample the value at posedge clk)";5�_�  �             �   f        ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�?     �   e   f           5�_�  �                f        ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�A     �   f   j   n       �   f   h   m    5�_�                  h   
    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�J     �   g   i   p      
covergroup5�_�                 h       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�Y     �   g   i   p      covergroup cg_supply @5�_�                 h   #    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�a     �   g   i   p      #covergroup cg_supply @(posedge clk)5�_�                 h   #    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�b     �   h   k   q          �   h   j   p    5�_�                 h       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�u     �   h   j   s          �   h   j   r    5�_�                 i       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�~     �   h   i              bins dd5�_�                 h        ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�     �   h   j   s          �   h   j   r    5�_�    	             i       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   i   k   t          �   i   k   s    5�_�    
          	   i       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   i   k   u          �   i   k   t    5�_�  	            
   j   '    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   i   k   u      '    supply_cpt : coverpoint inf.supply 5�_�  
               j   (    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   i   k   u      )    supply_cpt : coverpoint inf.supply {}5�_�                 j   (    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   i   m   u      )    supply_cpt : coverpoint inf.supply {}5�_�                 m       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   l   m          	    bins 5�_�                 k        ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   k   m   v    �   k   l   v    5�_�                 l       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   k   m   w      	    bins 5�_�                 k       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   j   k              5�_�                 k       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   j   l   v              bins 5�_�                 k       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   j   l   v              bins supply =5�_�                 k       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   j   l   v              bins supply ={}5�_�                 k       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��    �   j   l   v              bins supply ={[0:1023]}5�_�                 k       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   j   l   v              bins supply ={[0:1023]}5�_�                 k       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   k   m   w          �   k   m   v    5�_�                 l   )    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�o     �   l   n   x              �   l   n   w    5�_�                 o        ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2�     �   n   o           5�_�                 o        ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   o   r   x       �   o   q   w    5�_�                 q       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   p   r   y      cg_supply cg_supply_inst = new5�_�                 q       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   p   r   y       cg_supply cg_supply_inst = new()5�_�                 )       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   (   *   y      Dcovergroup cg_btn_size_cross @(posedge clk);// sample at posedge clk5�_�                 )       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   (   *   y      5covergroup cg_@(posedge clk);// sample at posedge clk5�_�                 )       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   (   *   y      <covergroup cg_window @(posedge clk);// sample at posedge clk5�_�                  )       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   (   *   y      Ecovergroup cg_window_btn_size @(posedge clk);// sample at posedge clk5�_�    !              )       ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   (   *   y      ?covergroup cg__btn_size @(posedge clk);// sample at posedge clk5�_�     "          !   q        ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   q   s   z       �   q   s   y    5�_�  !  #          "   r   7    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��     �   q   s   z      7cg_btn_size_led_ratio  cg_btn_size_led_ratio_inst = new5�_�  "  %          #   r   8    ����                                                                                                                =                                                                                                                                                                                                          d          d          V       Z2��    �   q   s   z      9cg_btn_size_led_ratio  cg_btn_size_led_ratio_inst = new()5�_�  #  &  $      %   r        ����                                                                                                                =                                                                                                                                                                                                          v           x           V        Z4w|     �   r   t   {       �   r   t   z    5�_�  %  '          &   s        ����                                                                                                                =                                                                                                                                                                                                          w           y           V        Z4w�     �   r   s          	cg_supply5�_�  &  (          '   v        ����                                                                                                                =                                                                                                                                                                                                          v           x           V        Z4w�     �   u   v          1cg_btn_size_cross cg_btn_size_cross_inst = new();   :cg_led            cg_led_inst            = new();            1cg_ratio_tran     cg_ratio_tran_inst     = new();5�_�  '  )          (   q       ����                                                                                                                =                                                                                                                                                                                                          v           v           V        Z4w�     �   p   r   w      !cg_supply cg_supply_inst = new();5�_�  (  *          )   p        ����                                                                                                                =                                                                                                                                                                                                          v           v           V        Z4w�   	 �   o   q   w       5�_�  )  +          *   s        ����                                                                                                                =                                                                                                                                                                                                          v           v           V        Z4x�     �   s   v   x       �   s   u   w    5�_�  *  ,          +   u       ����                                                                                                                =                                                                                                                                                                                                          x           x           V        Z4x�     �   s   u   y      4// ######################################### CHECKER   (########################################�   t   v   y      +// ########################################5�_�  +  -          ,   t   5    ����                                                                                                                =                                                                                                                                                                                                          w           w           V        Z4y     �   t   w   y      // �   t   v   x    5�_�  ,  .          -   v       ����                                                                                                                =                                                                                                                                                                                                          y           y           V        Z4y9     �   u   w   z      module Checker5�_�  -  /          .   v   *    ����                                                                                                                =                                                                                                                                                                                                          y           y           V        Z4yD     �   u   w   z      +module Checker(input clk, INF.CHECKER inf )5�_�  .  0          /   v   +    ����                                                                                                                =                                                                                                                                                                                                          y           y           V        Z4yE     �   u   w   z      +module Checker(input clk, INF.CHECKER inf )5�_�  /  1          0   v   +    ����                                                                                                                =                                                                                                                                                                                                          y           y           V        Z4yF     �   v   x   {       �   v   x   z    5�_�  0  2          1   v       ����                                                                                                                =                                                                                                                                                                                                          z           z           V        Z4yI     �   v   x   {    5�_�  1  3          2   w        ����                                                                                                                =                                                                                                                                                                                                          {           {           V        Z4y�     �   v   x   |       5�_�  2  4          3   w   J    ����                                                                                                                =                                                                                                                                                                                                          {           {           V        Z4y�     �   w   y   }          //�   w   y   |    5�_�  3  5          4   x       ����                                                                                                                =                                                                                                                                                                                                          |           |           V        Z4y�     �   w   y   }          property5�_�  4  6          5   x       ����                                                                                                                =                                                                                                                                                                                                          |           |           V        Z4y�     �   w   y   }          property()5�_�  5  7          6   x       ����                                                                                                                =                                                                                                                                                                                                          |           |           V        Z4y�     �   w   y   }          property()5�_�  6  8          7   x       ����                                                                                                                =                                                                                                                                                                                                          |           |           V        Z4y�   
 �   x   {   ~              �   x   z   }    5�_�  7  9          8   x       ����                                                                                                                =                                                                                                                                                                                                          ~           ~           V        Z4z     �   x   z   �              �   x   z       5�_�  8  :          9   y   	    ����                                                                                                                =                                                                                                                                                                                                                                V        Z4z     �   x   z   �      	        @5�_�  9  ;          :   y       ����                                                                                                                =                                                                                                                                                                                                                                V        Z4z$     �   x   z   �              @(posedge clk)5�_�  :  <          ;   y       ����                                                                                                                =                                                                                                                                                                                                                                V        Z4z$     �   x   z   �              @(posedge clk)5�_�  ;  =          <   y   #    ����                                                                                                                =                                                                                                                                                                                                                                V        Z4z)     �   x   z   �      #        @(posedge clk) inf.supply==5�_�  <  >          =   y   &    ����                                                                                                                =                                                                                                                                                                                                                                V        Z4z*     �   x   z   �      '        @(posedge clk) inf.supply=='d0'5�_�  =  ?          >   y   '    ����                                                                                                                =                                                                                                                                                                                                                                V        Z4z+     �   x   z   �      '        @(posedge clk) inf.supply=='d0'5�_�  >  @          ?   z        ����                                                                                                                =                                                                                                                                                                                                                                V        Z4{x     �   y   z           5�_�  ?  A          @   z       ����                                                                                                                =                                                                                                                                                                                                          ~           ~           V        Z4{y     �   z   |       5�_�  @  B          A   w       ����                                                                                                                =                                                                                                                                                                                                                                V        Z4{{     �   w   z   �          //�   w   y   �    5�_�  A  C          B   x       ����                                                                                                                =                                                                                                                                                                                                          �           �           V        Z4{     �   w   {   �          5�_�  B  D          C   y        ����                                                                                                                =                                                                                                                                                                                                          �           �           V        Z4{�     �   x   z   �       5�_�  C  E          D   y       ����                                                                                                                =                                                                                                                                                                                                          �           �           V        Z4{�     �   x   z   �              5�_�  D  F          E   y       ����                                                                                                                =                                                                                                                                                                                                          �           �           V        Z4{�     �   x   z   �              (inf.supply != 0)5�_�  E  G          F   y       ����                                                                                                                =                                                                                                                                                                                                          �           �           V        Z4{�    �   x   z   �              (inf.supply != 0)5�_�  F  H          G   }   '    ����                                                                                                                =                                                                                                                                                                                                          �           �           V        Z4|�     �   |   ~   �      '        @(posedge clk) inf.select_i != 5�_�  G  I          H   x        ����                                                                                                                =                                                                                                                                                                                                          x          z          V   *    Z4}9     �   w   x              sequence supply_seq;           (inf.supply != 0);       endsequence5�_�  H  J          I   {        ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}G     �   |   ~   �          supply_no_zero�   {   ~   �          �   {   }   �    5�_�  I  K          J   }       ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}m     �   |   ~   �          supply_no_zero5�_�  J  L          K   }       ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}t     �   |   ~   �          select_then_supply_no_zero5�_�  K  M          L   }   0    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}y     �   |   ~   �      0    select_then_supply_no_zero : assert property5�_�  L  N          M   }   6    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}}     �   |   ~   �      7    select_then_supply_no_zero : assert property(spec1)5�_�  M  O          N   }   7    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}     �   |      �      7    select_then_supply_no_zero : assert property(spec1)5�_�  N  P          O   ~   *    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   ~   �   �      %                                     �   ~   �   �    5�_�  O  Q          P           ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   ~   �   �       5�_�  P  R          Q      ,    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   ~   �   �      ,                                    $display5�_�  Q  S          R      -    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   ~   �   �      .                                    $display()5�_�  R  T          S      /    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   ~   �   �      0                                    $display("")5�_�  S  U          T      .    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   ~   �   �      0                                    $display("")5�_�  T  V          U      ?    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   ~   �   �      ?                                    $display("Spec_1 is wrong")5�_�  U  W          V   �   #    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4}�     �   �   �   �      !                                 �   �   �   �    5�_�  V  X          W      $    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4~     �      �   �      $                                    �      �   �    5�_�  W  Y          X   �   *    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4~
     �      �   �      *                                    $error5�_�  X  Z          Y   �   +    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4~     �      �   �      ,                                    $error()5�_�  Y  [          Z   �   -    ����                                                                                                                =                                                                                                                                                                                                          x          x          V   *    Z4~     �      �   �      .                                    $error("")5�_�  Z  \          [   �   +    ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~     �      �   �      .                                    $error("")   $                                 end�   �   �   �    5�_�  [  ]          \   �   =    ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~     �      �   �      =                                    $error("Spec_1 is wrong")5�_�  \  ^          ]      $    ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~    �   ~             @                                    $display("Spec_1 is wrong");5�_�  ]  _          ^   �       ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~:     �   �   �   �          //spec2. 5�_�  ^  `          _   �       ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~C     �   �   �   �      %    //changed from no_size_inf to any5�_�  _  a          `   �       ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~D     �   �   �   �      J    //spec2. When flavor_btn is not no_coffee, the required_size should be   #    changed from no_size_inf to any5�_�  `  b          a   �       ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~G     �   �   �   �      j    //spec2. When flavor_btn is not no_coffee, the required_size should be changed from no_size_inf to any       //other size requirement.5�_�  a  c          b   �   k    ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~H     �   �   �   �      �    //spec2. When flavor_btn is not no_coffee, the required_size should be changed from no_size_inf to any //other size requirement.5�_�  b  d          c   �   k    ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~I     �   �   �   �          //�   �   �   �    5�_�  c  e          d   ~   &    ����                                                                                                                =                                                                                                                                                                                                             .          <          <    Z4~j     �   ~   �   �      %                                     �   ~   �   �    5�_�  d  f          e      *    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~q     �   ~   �   �      *                                    $error5�_�  e  g          f      +    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~s     �   ~   �   �      ,                                    $error()5�_�  f  h          g      -    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~s     �   ~   �   �      .                                    $error("")5�_�  g  i          h      ,    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~t     �   ~   �   �      .                                    $error("")5�_�  h  j          i   �   =    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~w     �      �   �      =                                    other size requirement.")5�_�  i  k          j      %    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~z     �   ~   �   �      �                                    $error("When flavor_btn is not no_coffee, the required_size should be changed from no_size_inf to any5�_�  j  l          k   �   %    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   �   �   �      >                                    $error("Spec_1 is wrong");5�_�  k  m          l      %    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   ~   �   �      �                                    $display("When flavor_btn is not no_coffee, the required_size should be changed from no_size_inf to any5�_�  l  n          m   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   �   �          @                                    $display("Spec_1 is wrong");5�_�  m  o          n   ~   !    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   ~   �   �    �   ~      �    5�_�  n  p          o   �        ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   �   �   �       5�_�  o  q          p   �   	    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   �   �   �      	        @5�_�  p  s          q   �   
    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   �   �   �              @()5�_�  q  t  r      s   �   
    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   �   �   �              @()5�_�  s  u          t   �       ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   �   �   �              @(posedge clk)5�_�  t  v          u   �   3    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4    �   �   �   �      3        @(posedge clk) inf.flavor_btn != no_coffee 5�_�  u  w          v   �       ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4y     �   �   �   �          flavor_btn_ required_size�   �   �   �          �   �   �   �    5�_�  v  x          w   �       ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �          flavor_btn_ required_size5�_�  w  y          x   �       ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �          flavor_btn_ required_size5�_�  x  z          y   �   !    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �      !    flavor_btn_then_required_size5�_�  y  {          z   �   3    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �      3    flavor_btn_then_required_size : assert property5�_�  z  |          {   �   9    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �      :    flavor_btn_then_required_size : assert property(spec2)5�_�  {  }          |   �   9    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �          �   �   �   �    5�_�  |  ~          }   �   -    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �      (                                        �   �   �   �    5�_�  }            ~   �   &    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4�     �   �   �   �    5�_�  ~  �             �        ����                                                                                                                =                                                                                                                                                                                                             (       �   $       V   (    Z4�     �   �   �   �    �   �   �   �    5�_�    �          �   �   3    ����                                                                                                                =                                                                                                                                                                                                             (       �   $       V   (    Z4�     �   �   �   �      @                                    $display("Spec_1 is wrong");5�_�  �  �          �   �   ,    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   -          -    Z4�     �   �   �   �      �                                    $error("When flavor_btn is not no_coffee, the required_size should be changed from no_size_inf to any5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   -          -    Z4�     �   �   �   �      ,                                    $error("   >                                    other size requirement.");5�_�  �  �          �   �   ,    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      G                                    $error(" other size requirement.");5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      /                                    $error("");�   �   �   �    5�_�  �  �          �   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �          '                                    end5�_�  �  �          �   �   "    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      $                                 end5�_�  �  �          �   �   !    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�    �   �   �   �      $                                 end5�_�  �  �          �   �   #    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      $                                    �   �   �   �    5�_�  �  �          �   �   &    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      E    //spec3. The next flavor_btn or select_i should be inserted after   '    //out_valid is low within 1~3 cycle5�_�  �  �          �   �   F    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      i    //spec3. The next flavor_btn or select_i should be inserted after //out_valid is low within 1~3 cycle5�_�  �  �          �   �   E    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �          //�   �   �   �    5�_�  �  �          �   �   !    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�!     �   �   �   �      !    out_valid_1to3_then_select_i:5�_�  �  �          �   �   !    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�$     �   �   �   �          //�   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�+     �   �   �   �              �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�.     �   �   �   �              �   �   �   �    5�_�  �  �          �   �   	    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�0     �   �   �   �      	        @5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�2     �   �   �   �              @(posedge)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�3     �   �   �   �              @(posedge)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�5     �   �   �   �              @(posedge clk)5�_�  �  �          �   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�p     �   �   �   �      )        @(posedge clk) inf.out_valid |=> 5�_�  �  �          �   �   .    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      .        @(posedge clk) inf.out_valid == 0 |=> 5�_�  �  �          �   �   /    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      0        @(posedge clk) inf.out_valid == 0 |=> []5�_�  �  �          �   �   /    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      0        @(posedge clk) inf.out_valid == 0 |=> []5�_�  �  �          �   �   2    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      3        @(posedge clk) inf.out_valid == 0 |=> [1:3]5�_�  �  �          �   �   0    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      3        @(posedge clk) inf.out_valid == 0 |=> [1:3]5�_�  �  �          �   �   .    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      3        @(posedge clk) inf.out_valid == 0 |=> [1:3]5�_�  �  �          �   �   .    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      5        @(posedge clk) inf.out_valid == 0 |=> ##[1:3]5�_�  �  �          �   �   3    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      6        @(posedge clk) inf.out_valid == 0 |=> (##[1:3]5�_�  �  �          �   �   5    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      6        @(posedge clk) inf.out_valid == 0 |=> (##[1:3]5�_�  �  �          �   �   6    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      6        @(posedge clk) inf.out_valid == 0 |=> (##[1:3]5�_�  �  �          �   �   6    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      8        @(posedge clk) inf.out_valid == 0 |=> (##[1:3] )5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �          endproperty5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �          endproperty5�_�  �  �          �   {       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   z   |   �          endproperty5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�"     �   �   �   �          endproperty: spe35�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �              �   �   �   �    5�_�  �  �          �   �   7    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      S        @(posedge clk) inf.out_valid == 0 |=> (##[1:3] flavor_btn or inf.select_i )5�_�  �  �          �   �   7    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      S        @(posedge clk) inf.out_valid == 0 |=> (##[1:3] flavor_btn or inf.select_i )5�_�  �  �          �   �   R    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      T        @(posedge clk) inf.out_valid == 0 |=> (##[1:3] (flavor_btn or inf.select_i )5�_�  �  �          �   �   S    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      S        @(posedge clk) inf.out_valid == 0 |=> (##[1:3] (flavor_btn or inf.select_i)5�_�  �  �          �   �   U    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      U        @(posedge clk) inf.out_valid == 0 |=> (##[1:3] (flavor_btn or inf.select_i) )5�_�  �  �          �   �   !    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �    5�_�  �  �          �   �   "    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      "    out_valid_1to3_then_select_i: 5�_�  �  �          �   �   1    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      1    out_valid_1to3_then_select_i: assert property5�_�  �  �          �   �   7    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      8    out_valid_1to3_then_select_i: assert property(spec3)5�_�  �  �          �   �   8    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      8    out_valid_1to3_then_select_i: assert property(spec3)5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �       5�_�  �  �          �   �   ,    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      ,                                    $display5�_�  �  �          �   �   -    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      .                                    $display()5�_�  �  �          �   �   /    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      0                                    $display("")5�_�  �  �          �   �   .    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      0                                    $display("")5�_�  �  �          �   �   >    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      >                                    $display("Spec3 is wrong")5�_�  �  �          �   �   >    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      $                                    �   �   �   �    5�_�  �  �          �   �   *    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      *                                    $error5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      ,                                    $error()5�_�  �  �          �   �   -    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      .                                    $error("")5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      .                                    $error("")�   �   �   �    5�_�  �  �          �   �   �    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      �                                    $error("The next flavor_btn or select_i should be inserted after out_valid is low within 1~3 cycle")5�_�  �  �          �   �   �    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      $                                    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��    �   �   �   �      #                                end5�_�  �  �  �      �   �   	    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      	endmodule5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �          
endmodule:5�_�  �  �          �   v        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�$     �   u   v          ,module Checker(input clk, INF.CHECKER inf );5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�E     �   �   �   �      "                                  �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�R     �   �   �   �          endproperty5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�[     �   �   �   �       5�_�  �  �          �   �   	    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�^     �   �   �   �      	        @5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�l     �   �   �   �       5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�s     �   �   �   �      @    //After rst_n signal, all output should be zero immediately.5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�y     �   �   �   �              @(posedge clk)5�_�  �  �          �   �   
    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �              @(posedge clk) rst_n5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �              @(negedge clk) rst_n5�_�  �  �          �   �   "    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      "        @(negedge inf.rst_n) rst_n5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�0     �   �   �   �              @(negedge inf.rst_n) 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�4     �   �   �   �              @(negedge inf.rst_n) 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�E     �   �   �   �              inf.out_valid == 0) 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�E     �   �   �   �              inf.out_valid == 0) 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�G     �   �   �   �              inf.out_valid == 0) 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�L     �   �   �   �              (inf.out_valid == 0) 5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�R     �   �   �   �               (inf.out_valid == 0) or 5�_�  �  �          �   �   !    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�R     �   �   �   �      "        (inf.out_valid == 0) or ()5�_�  �  �          �   �   !    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�T     �   �   �   �      "        (inf.out_valid == 0) or ()5�_�  �  �          �   �   %    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�e     �   �   �   �      2        (inf.out_valid == 0) or (inf.flavor_btn==)5�_�  �  �          �   �   1    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�i     �   �   �   �      2        (inf.out_valid == 0) or (inf.flavor_out==)5�_�  �  �          �   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�m     �   �   �   �      ;        (inf.out_valid == 0) or (inf.flavor_out==no_coffee)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      <        (inf.out_valid == 0) or (inf.flavor_out==no_coffee) 5�_�  �  �          �   �   =    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      =        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) 5�_�  �  �          �   �   A    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      A        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and 5�_�  �  �          �   �   B    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      C        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and ()5�_�  �  �          �   �   B    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      C        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and ()5�_�  �  �          �   �   Q    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      R        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and (inf.select_i ==)5�_�  �  �          �   �   B    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      C        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and ()5�_�  �  �          �   �   @    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      @        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and5�_�  �  �          �   �   A    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      A        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and 5�_�  �  �          �   �   B    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      C        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and ()5�_�  �  �          �   �   A    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      C        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and ()5�_�  �  �          �   �   	    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      
        ()5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      A        (inf.out_valid == 0) and (inf.flavor_out==no_coffee) and 5�_�  �  �          �   �   3    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      B        (inf.out_valid === 0) and (inf.flavor_out==no_coffee) and 5�_�  �  �          �   �   &    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      V        @(posedge clk) inf.out_valid == 0 |=> (##[1:3] (flavor_btn or inf.select_i) );5�_�  �  �          �   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      %        (inf.window.espresso.led ===)5�_�  �  �          �   �   M    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      M        (inf.window.espresso.led === red && inf.window.espresso.monitor == 0)5�_�  �  �          �   �   P    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4��     �   �   �   �      Q        (inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and5�_�  �  �          �   �   3    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      M        (inf.window.milk.led === red && inf.window.espresso.monitor == 0) and5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      Q        (inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and5�_�  �  �          �   �   8    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      R        (inf.window.chocolate.led === red && inf.window.espresso.monitor == 0) and5�_�  �  �          �   �   7    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      Q        (inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �   �      N        (inf.window.espresso.led === red && inf.window.froth.monitor == 0) and5�_�  �  �          �   �   K    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�&     �   �   �   �      K        (inf.window.froth.led === red && inf.window.froth.monitor == 0) and5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�7     �   �   �   �          �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�S     �   �   �   �           rst_n_check: assert property5�_�  �  �          �   �   &    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�V     �   �   �   �      '    rst_n_check: assert property(spec4)5�_�  �  �          �   �   &    ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�W     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�\     �   �   �   �                           �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�]     �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�b     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�h     �   �   �   �      ?                                    $display("Spec3 is wrong");5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�h     �   �   �   �      �                                    $error("The next flavor_btn or select_i should be inserted after out_valid is low within 1~3 cycle");5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�i     �   �   �           5�_�  �  �          �   �   $    ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�l     �   �   �   �      1                      $display("Spec3 is wrong");5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�o     �   �   �   �      {                      $error("The next flavor_btn or select_i should be inserted after out_valid is low within 1~3 cycle");5�_�  �             �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�x     �   �   �   �      !                      $error("");�   �   �   �    5�_�  �                �   0    ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4��     �   �   �   �    5�_�                  �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4��     �   �   �   �    �   �   �   �    5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      Q        (inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and   I        (inf.window.milk.led === red && inf.window.milk.monitor == 0) and   S        (inf.window.chocolate.led === red && inf.window.chocolate.monitor == 0) and   H        (inf.window.froth.led === red && inf.window.froth.monitor == 0);�   �   �   �      C        (inf.out_valid === 0) and (inf.flavor_out===no_coffee) and 5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      S                        (inf.out_valid === 0) and (inf.flavor_out===no_coffee) and 5�_�                 �   4    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      U                        if(inf.out_valid === 0) and (inf.flavor_out===no_coffee) and 5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �    5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      a                        (inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and5�_�    	             �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      d                        if (inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and5�_�    
        	   �   7    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      ;                        if(inf.flavor_out===no_coffee) and 5�_�  	            
   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �    5�_�  
               �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                                  �   �   �   �    5�_�                 �   $    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      $                            $display5�_�                 �   %    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      &                            $display()5�_�                 �   )    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      /                        if(inf.out_valid === 0)5�_�                 �   %    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      &                            $display()5�_�                 �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �    �   �   �   �    5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      1                      $display("Spec4 is wrong");�   �   �   �    5�_�                 �   \    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      n                      $display("After rst_n signal, all output should be zero immediately.");Spec4 is wrong");5�_�                 �   \    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      \                      $display("After rst_n signal, all output should be zero immediately.")5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �          [                      $error("After rst_n signal, all output should be zero immediately.");5�_�                 �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �           5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �                              �   �   �   �    5�_�                 �   %    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      &                            $display()5�_�                 �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      (                            $display("")5�_�                 �   4    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      5                            $display("out_valid: %d")5�_�                 �   C    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�"     �   �   �   �      C                            $display("out_valid: %d",inf.out_valid)5�_�                 �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�#     �   �   �           5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�&     �   �   �   �    �   �   �   �    5�_�                 �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�(     �   �   �   �      D                            $display("out_valid: %d",inf.out_valid);5�_�                 �   :    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�.     �   �   �   �      E                            $display("flavor_out: %d",inf.out_valid);5�_�                  �   )    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�5     �   �   �   �      6                        if(inf.flavor_out===no_coffee)5�_�    !              �   +    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�6     �   �   �   �      7                        if(inf.flavor_out ===no_coffee)5�_�     "          !   �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�:     �   �   �           5�_�  !  #          "   �   3    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�=     �   �   �   �      c                        if(inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and5�_�  "  $          #   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�@     �   �   �   �      c                        if(inf.window.espresso.led !== red && inf.window.espresso.monitor == 0) and5�_�  #  %          $   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�D     �   �   �   �                                  5�_�  $  &          %   �   $    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�F     �   �   �   �      $                            $display5�_�  %  '          &   �   %    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�F     �   �   �   �      &                            $display()5�_�  &  (          '   �   %    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�H     �   �   �   �      &                            $display()5�_�  '  )          (   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�N     �   �   �   �      (                            $display("")5�_�  (  *          )   �   7    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�^     �   �   �   �      8                            $display("espresso.led: %s")5�_�  )  +          *   �   P    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�n     �   �   �   �      P                            $display("espresso.led: %s",inf.window.espresso.led)5�_�  *  ,          +   �   P    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�o     �   �   �   �                              �   �   �   �    5�_�  +  -          ,   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�s     �   �   �   �                              if   D                            && inf.window.espresso.monitor == 0) and5�_�  ,  .          -   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�t     �   �   �   �      C                        if && inf.window.espresso.monitor == 0) and5�_�  -  /          .   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�u     �   �   �   �      @                        if inf.window.espresso.monitor == 0) and5�_�  .  0          /   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�u     �   �   �   �      @                        if inf.window.espresso.monitor == 0) and5�_�  /  1          0   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�v     �   �   �   �      @                        if inf.window.espresso.monitor == 0) and5�_�  0  2          1   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�w     �   �   �   �      B                        if() inf.window.espresso.monitor == 0) and5�_�  1  3          2   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�w     �   �   �   �      B                        if() inf.window.espresso.monitor == 0) and5�_�  2  4          3   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�x     �   �   �   �      A                        if( inf.window.espresso.monitor == 0) and5�_�  3  5          4   �   >    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�|     �   �   �   �      @                        if(inf.window.espresso.monitor == 0) and5�_�  4  6          5   �   =    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�|     �   �   �   �      >                        if(inf.window.espresso.monitor == 0) a5�_�  5  7          6   �   <    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�}     �   �   �   �    5�_�  6  8          7   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �    �   �   �   �    5�_�  7  9          8   �   /    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      Q                            $display("espresso.led: %s",inf.window.espresso.led);5�_�  8  :          9   �   P    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      U                            $display("espresso.monitor: %s",inf.window.espresso.led);5�_�  9  ;          :   �   9    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      Y                            $display("espresso.monitor: %s",inf.window.espresso.monitor);5�_�  :  <          ;   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      Y                        (inf.window.milk.led === red && inf.window.milk.monitor == 0) and5�_�  ;  =          <   �   6    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      [                        if(inf.window.milk.led === red && inf.window.milk.monitor == 0) and5�_�  <  >          =   �   /    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      \                        if(inf.window.milk.led === red) && inf.window.milk.monitor == 0) and5�_�  =  ?          >   �   6    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      =                        if(inf.window.espresso.monitor == 0) 5�_�  >  @          ?   �   6    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      >                        if(inf.window.espresso.monitor! == 0) 5�_�  ?  A          @   �   9    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      ?                        if(inf.window.espresso.monitor ! == 0) 5�_�  @  B          A   �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �           5�_�  A  C          B   �   8    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      \                        if(inf.window.milk.led !== red) && inf.window.milk.monitor == 0) and5�_�  B  D          C   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                                  5�_�  C  E          D   �   $    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      $                            $display5�_�  D  F          E   �   %    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      &                            $display()5�_�  E  G          F   �   %    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      &                            $display()5�_�  F  H          G   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      (                            $display("")5�_�  G  I          H   �   .    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      0                            $display("milk.led")5�_�  H  J          I   �   3    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      4                            $display("milk.led: %s")5�_�  I  K          J   �   H    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      H                            $display("milk.led: %s",inf.window.milk.led)5�_�  J  L          K   �   H    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                              �   �   �   �    5�_�  K  M          L   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                              if   @                            && inf.window.milk.monitor == 0) and5�_�  L  N          M   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      ?                        if && inf.window.milk.monitor == 0) and5�_�  M  O          N   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      <                        if inf.window.milk.monitor == 0) and5�_�  N  P          O   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      <                        if inf.window.milk.monitor == 0) and5�_�  O  Q          P   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      =                        if (inf.window.milk.monitor == 0) and5�_�  P  R          Q   �   <    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      <                        if(inf.window.milk.monitor == 0) and5�_�  Q  S          R   �   3    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      8                        if(inf.window.milk.monitor == 0)5�_�  R  T          S   �   4    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      8                        if(inf.window.milk.monitor != 0)5�_�  S  U          T   �   4    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �    �   �   �   �    5�_�  T  V          U   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      Y                            $display("espresso.monitor: %d",inf.window.espresso.monitor);5�_�  U  W          V   �   C    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      U                            $display("milk.monitor: %d",inf.window.espresso.monitor);5�_�  V  X          W   �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �           5�_�  W  Y          X   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      c                        (inf.window.chocolate.led === red && inf.window.chocolate.monitor == 0) and5�_�  X  Z          Y   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�      �   �   �   �      e                        if(inf.window.chocolate.led === red && inf.window.chocolate.monitor == 0) and5�_�  Y  [          Z   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �    �   �   �   �    5�_�  Z  \          [   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�	     �   �   �   �      I                            $display("milk.led: %s",inf.window.milk.led);5�_�  [  ]          \   �   4    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      <                        if(inf.window.chocolate.led === red)5�_�  \  ^          ]   �   D    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      N                            $display("chocolate.led: %s",inf.window.milk.led);5�_�  ]  _          ^   �   L    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �                              �   �   �   �    5�_�  ^  `          _   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �                              if5�_�  _  a          `   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �                              if()5�_�  `  b          a   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �                              if()5�_�  a  c          b   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �                              if(                              5�_�  b  d          c   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �                              if(    E                            && inf.window.chocolate.monitor == 0) and5�_�  c  e          d   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�      �   �   �   �      E                        if( && inf.window.chocolate.monitor == 0) and5�_�  d  f          e   �   9    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�$     �   �   �   �      B                        if( inf.window.chocolate.monitor == 0) and5�_�  e  g          f   �   >    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�$     �   �   �   �      C                        if( inf.window.chocolate.monitor !== 0) and5�_�  f  h          g   �   ?    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�%     �   �   �   �      C                        if( inf.window.chocolate.monitor !== 0) and5�_�  g  i          h   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�'     �   �   �   �      ?                        if( inf.window.chocolate.monitor !== 0)5�_�  h  k          i   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�,     �   �   �   �    �   �   �   �    5�_�  i  l  j      k   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�5     �   �   �   �      Q                            $display("milk.monitor: %d",inf.window.milk.monitor);5�_�  k  m          l   �   H    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�9     �   �   �   �      V                            $display("chocolate.monitor: %d",inf.window.milk.monitor);5�_�  l  n          m   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�=     �   �   �   �      <                        if(inf.window.chocolate.led !== red)5�_�  m  o          n   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�@     �   �   �                                      and5�_�  n  p          o   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�E     �   �   �   �    �   �   �   �    5�_�  o  q          p   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�F     �   �   �   �      S                            $display("chocolate.led: %s",inf.window.chocolate.led);5�_�  p  r          q   �   @    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�I     �   �   �   �      O                            $display("froth.led: %s",inf.window.chocolate.led);5�_�  q  s          r   �   D    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�K     �   �   �   �                              �   �   �   �    5�_�  r  t          s   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�M     �   �   �   �                              if5�_�  s  u          t   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�O     �   �   �   �                              if()5�_�  t  v          u   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�P     �   �   �                                  if()5�_�  u  w          v   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�Q     �   �   �   �      X                        (inf.window.froth.led === red && inf.window.froth.monitor == 0);5�_�  v  x          w   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�[     �   �   �   �      Z                        if(inf.window.froth.led === red && inf.window.froth.monitor == 0);5�_�  w  y          x   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�\     �   �   �   �      =                        if(&& inf.window.froth.monitor == 0);5�_�  x  z          y   �   :    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�_     �   �   �   �      :                        if(inf.window.froth.monitor == 0);5�_�  y  {          z   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�c     �   �   �   �    �   �   �   �    5�_�  z  |          {   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�d     �   �   �   �      [                            $display("chocolate.monitor: %d",inf.window.chocolate.monitor);5�_�  {  }          |   �   D    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�h     �   �   �   �      W                            $display("froth.monitor: %d",inf.window.chocolate.monitor);5�_�  |  ~          }   �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�l     �   �   �           5�_�  }            ~   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�}     �   �   �                              $fatal;5�_�  ~  �             �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                       �   �   �   �    5�_�    �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �              �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      //  spec5 After flavor_btn 5�_�  �  �          �   �   F    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      F//  spec5 After flavor_btn (also depends on ratio signal) or select_i 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      //  last one)5�_�  �  �          �   �   
    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      J//  spec5 After flavor_btn (also depends on ratio signal) or select_i (the5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �              �   �   �   �    5�_�  �  �          �   �   	    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      	        @5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �              @(posedge clk)5�_�  �  �          �   �   &    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�H     �   �   �   �      &        @(posedge clk) inf.flavor_btn 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�U     �   �   �   �      4        @(posedge clk) inf.flavor_btn !== no_coffee)5�_�  �  �          �   �   5    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�\     �   �   �   �      5        @(posedge clk) (inf.flavor_btn !== no_coffee)5�_�  �  �          �   �   :    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�`     �   �   �   �      :        @(posedge clk) (inf.flavor_btn !== no_coffee) and 5�_�  �  �          �   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�`     �   �   �   �      <        @(posedge clk) (inf.flavor_btn !== no_coffee) and ()5�_�  �  �          �   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�f     �   �   �   �      <        @(posedge clk) (inf.flavor_btn !== no_coffee) and ()5�_�  �  �          �   �   D    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�o     �   �   �   �      E        @(posedge clk) (inf.flavor_btn !== no_coffee) and (select_i )5�_�  �  �          �   �   H    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      I        @(posedge clk) (inf.flavor_btn !== no_coffee) and (select_i !== )5�_�  �  �          �   �   M    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      M        @(posedge clk) (inf.flavor_btn !== no_coffee) and (select_i !== none)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      N        @(posedge clk) (inf.flavor_btn !== no_coffee) and (select_i !== none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      P        @(posedge clk) ()(inf.flavor_btn !== no_coffee) and (select_i !== none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      P        @(posedge clk) ()(inf.flavor_btn !== no_coffee) and (select_i !== none))5�_�  �  �          �   �   O    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      O        @(posedge clk) ((inf.flavor_btn !== no_coffee) and (select_i !== none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                             �   �   �   �    5�_�  �  �          �   �   (    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      R        @(posedge clk) ((inf.flavor_btn !== no_coffee) and (select_i !== none)) or5�_�  �  �          �   �   E    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      R                       ((inf.flavor_btn !== no_coffee) and (select_i !== none)) or5�_�  �  �          �   �   R    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      R                       ((inf.flavor_btn !== no_coffee) and (select_i === none)) or5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      R        @(posedge clk) ((inf.flavor_btn === no_coffee) and (select_i !== none)) or5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      T        @(posedge clk)() ((inf.flavor_btn === no_coffee) and (select_i !== none)) or5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      T        @(posedge clk)() ((inf.flavor_btn === no_coffee) and (select_i !== none)) or5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      S        @(posedge clk)( ((inf.flavor_btn === no_coffee) and (select_i !== none)) or5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �           5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                         )5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                         ) |=> 5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                         ) |=> ()5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                         ) |=> ()5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                         ) |=> (##)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                         ) |=> (##[])5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                         ) |=> (##[])5�_�  �  �          �   �   "    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      #                   ) |=> (##[1:30])5�_�  �  �          �   �   -    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      -                   ) |=> (##[1:30] out_valid)5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �           5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      .                   ) |=> (##[1:30] out_valid);5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      R                       ((inf.flavor_btn === no_coffee) and (select_i !== none)) or5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      O                       ((inf.flavor_btn !== no_coffee) and (select_i === none))5�_�  �  �          �   �   J    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      J                       ((inf.flavor_btn !== none) and (select_i === none))5�_�  �  �          �   �   L    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      M                       ((inf.flavor_btn !== none) and (select_i === none)) or5�_�  �  �          �   �   K    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�      �   �   �   �                             5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�      �   �   �   �                             ()5�_�  �  �          �   �   2    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      3                       ((inf.flavor_btn === ratio))5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      7                       ((inf.flavor_btn === ratio) and)5�_�  �  �          �   �   <    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      =                       ((inf.flavor_btn === user_define) and)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �          >                       ((inf.flavor_btn === user_define) and )5�_�  �  �          �   �   '    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      M                       ((inf.flavor_btn === none) and (select_i !== none)) or5�_�  �  �          �   �   0    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      M                       ((inf.flavor_btn === none) and (select_i !== none)) or5�_�  �  �          �   �   0    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      M                       ((inf.flavor_btn === none) and (select_i !== none)) or5�_�  �  �          �   �   0    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      M                       ((inf.flavor_btn !== none) and (select_i === none)) or5�_�  �  �          �   �   p    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      p                       ((inf.flavor_btn !== none && inf.flavor_btn !== user_define ) and (select_i === none)) or5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �          property spec5;5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4��     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�     �   �   �   �      )    property spec5_supply_general_coffee;5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�     �   �   �   �          property spec5_5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�     �   �   �   �          endproperty5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�     �   �   �   �      +    endproperty spec5_supply_general_coffee5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�     �   �   �          M                       ((inf.flavor_btn === none) and (select_i !== none)) or5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�"     �   �   �   �      m                       ((inf.flavor_btn !== none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�#     �   �   �   �      j                       ((.flavor_btn !== none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�#     �   �   �   �      i                       ((flavor_btn !== none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�$     �   �   �   �      ^                       ((!== none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�%     �   �   �   �      Z                       ((none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�%     �   �   �   �      U                       ((&& inf.flavor_btn !== user_define ) and (select_i === none))5�_�  �  �          �   �   (    ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�+     �   �   �   �      R                       ((inf.flavor_btn !== user_define ) and (select_i === none))5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�<     �   �   �   �      .                   ) |=> (##[0:30] out_valid);5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�?     �   �   �   �      .                   ) |=> (##[4:30] out_valid);5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�A     �   �   �   �      .                   ) |=> (##[4:34] out_valid);5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�C     �   �   �   �      .                   ) |=> (##[3:34] out_valid);5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�\     �   �   �   �      .                   ) |=> (##[3:33] out_valid);5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�]     �   �   �   �      .                   ) |=> (##[3:34] out_valid);5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�_     �   �   �   �      .                   ) |=> (##[3:33] out_valid);5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�t     �   �   �   �          �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�~     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4��     �   �   �   �          out_valid_cycle_check:5�_�  �  �          �   �   *    ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4��     �   �   �   �      *    out_valid_cycle_check: assert property5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4��     �   �   �   �      ,    out_valid_cycle_check: assert property()5�_�  �  �          �   �   +    ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4��     �   �   �   �      ,    out_valid_cycle_check: assert property()5�_�  �  �          �   �   G    ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�     �   �   �   �      G    out_valid_cycle_check: assert property(spec5_supply_general_coffee)5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      ]                      $display("After rst_n signal, all output should be zero immediately.");�   �   �   �      1                      $display("Spec4 is wrong");5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �           5�_�  �  �          �   �   .    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�     �   �   �   �      ;                                $display("Spec4 is wrong");5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �   .       �          V   .    Z4�&     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �                 Z4�.     �   �   �   �      D//  After flavor_btn (also depends on ratio signal) or select_i (the   $//  last one) is high, the out_valid   //  should be high in 30 cycle.5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �                 Z4�0     �   �   �   �      @After flavor_btn (also depends on ratio signal) or select_i (the5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �                 Z4�1     �   �   �   �       last one) is high, the out_valid�   �   �   �      @After flavor_btn (also depends on ratio signal) or select_i (the5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �                 Z4�4     �   �   �   �      should be high in 30 cycle.5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �                 Z4�7     �   �   �   �      A"After flavor_btn (also depends on ratio signal) or select_i (the    last one) is high, the out_valid5�_�  �  �          �   �   A    ����                                                                                                                =                                                                                                                                                                                                          �           �                 Z4�8     �   �   �   �      b"After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid   should be high in 30 cycle."5�_�  �  �          �   �   d    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�A     �   �   �   �      g                                $display("After rst_n signal, all output should be zero immediately.");5�_�  �  �          �   �   )    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�E     �   �   �   �      f                                $display("After rst_n signal, all output should be zero immediately.);5�_�  �  �  �      �   �   (    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�V     �   �   �   �    �   �   �   �    5�_�  �  �          �   �   )    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�Z     �   �   �   �      +                                $display();5�_�  �  �          �   �   (    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�[     �   �   �   �       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�^     �   �   �   �      "After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle."   );5�_�  �  �          �   �   (    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�_     �   �   �   �      )                                $display(   �"After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�b    �   �   �          "After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle."5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�g     �   �   �           5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�g     �   �   �           5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�h     �   �   �           5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�h     �   �   �           5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�}     �   �   �   �                                 �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4��     �   �   �   �      G    out_valid_cycle_check: assert property(spec5_supply_general_coffee)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4��     �   �   �   �          out_valid_cycle_check5�_�  �  �          �   �        ����                                                                                                                =                                                                                                                                                                                                          �           �          V        Z4��     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �          V        Z4��     �   �   �   �      ]    out_valid_cycle_check_general_coffee_supply: assert property(spec5_supply_general_coffee)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �          V        Z4��     �   �   �   �      2    : assert property(spec5_supply_general_coffee)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �           �          V        Z4��     �   �   �   �      !    out_valid_cycle_check_custom:   0    assert property(spec5_supply_general_coffee)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      ;                                $display("Spec5 is wrong");   �                                $display( "After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");�   �   �   �      %                           else begin5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                                 end5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �                                 end5�_�  �  �          �   �   2    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      N    out_valid_cycle_check_custom: assert property(spec5_supply_general_coffee)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      D    out_valid_cycle_check_custom: assert property(spec5_user_define)5�_�  �  �          �   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      >    out_valid_cycle_check_: assert property(spec5_user_define)5�_�  �  �          �   �   <    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                                $display( "After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�  �  �          �   �   <    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                                $display( "After flavor_btn ) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�  �            �   �   <    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                                $display( "After flavor_btn  or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�  �              �   D    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                                         $display( "After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�               �   R    ����                                                                                                                =                                                                                                                                                                                                          �   R       �   �          �    Z4��     �   �   �   �      �                                         $display( "After flavor_btn==user_define (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�                 �   Q    ����                                                                                                                =                                                                                                                                                                                                          �   R       �   �          �    Z4��    �   �   �   �      �                                         $display( "After flavor_btn==user_define  is high, the out_valid should be high in 30 cycle.");5�_�                 �   R    ����                                                                                                                =                                                                                                                                                                                                          �   R       �   X          X    Z4��     �   �   �   �      �                                         $display( "After flavor_btn==user_define is high, the out_valid should be high in 30 cycle.");5�_�    	             �   Q    ����                                                                                                                =                                                                                                                                                                                                          �   R       �   X          X    Z4�      �   �   �   �      �                                         $display( "After flavor_btn==user_define , the out_valid should be high in 30 cycle.");5�_�    
          	   �   R    ����                                                                                                                =                                                                                                                                                                                                          �   R       �   X          X    Z4�     �   �   �   �                                               $display( "After flavor_btn==user_define, the out_valid should be high in 30 cycle.");5�_�  	            
   �   (    ����                                                                                                                =                                                                                                                                                                                                          �   R       �   X          X    Z4�     �   �   �   �      ]    out_valid_cycle_check_general_coffee_supply: assert property(spec5_supply_general_coffee)5�_�  
             �   @    ����                                                                                                                =                                                                                                                                                                                                          �   @       �   F          F    Z4�     �   �   �   �      V    out_valid_cycle_check_general_coffee: assert property(spec5_supply_general_coffee)5�_�               �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�)     �   �   �   �      )    property spec5_supply_general_coffee;5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�6     �   �   �          M                       ((inf.flavor_btn === none) and (select_i !== none)) or5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�>     �   �   �   �      ,    endproperty :spec5_supply_general_coffee5�_�                 �        ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�B     �   �   �   �    �   �   �   �    5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�C     �   �   �   �    5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�H     �   �   �   �      "    property spec5_general_coffee;5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�H     �   �   �   �          property spec5_general_;5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�L     �   �   �   �      %    endproperty :spec5_general_coffee5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �          V       Z4�M     �   �   �   �          endproperty :spec5_general_5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�S     �   �   �   �      "    property spec5_general_supply;5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�T     �   �   �   �          property spec5__supply;5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�W     �   �   �   �      %    endproperty :spec5_general_supply5�_�                 �   (    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�d     �   �   �   �      m                       ((inf.flavor_btn !== none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�                 �   4    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�q     �   �   �   �      m                       ((inf.flavor_btn === none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�                 �   1    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�r     �   �   �   �      M                       ((inf.flavor_btn === none &&  and (select_i === none))5�_�                 �   1    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�s     �   �   �   �      L                       ((inf.flavor_btn === none &  and (select_i === none))5�_�                 �   1    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�s     �   �   �   �      K                       ((inf.flavor_btn === none   and (select_i === none))5�_�                  �   1    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�u     �   �   �   �      J                       ((inf.flavor_btn === none  and (select_i === none))5�_�    !              �   I    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      I                       ((inf.flavor_btn === none and (select_i === none))5�_�     "          !   �   ?    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      M                       ((inf.flavor_btn === none and (select_i === none)) |=>5�_�  !  #          "   �   M    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      M                       ((inf.flavor_btn === none and (select_i !== none)) |=>5�_�  "  $          #   �   Q    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      Q                       ((inf.flavor_btn === none and (select_i !== none)) |=> ###5�_�  #  %          $   �   U    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      V                       ((inf.flavor_btn === none and (select_i !== none)) |=> ###[0:3]5�_�  $  &          %   �   Q    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      V                       ((inf.flavor_btn === none and (select_i !== none)) |=> ###[0:3]5�_�  %  '          &   �   U    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      U                       ((inf.flavor_btn === none and (select_i !== none)) |=> ##[0:3]5�_�  &  (          '   �   N    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      h                       ((inf.flavor_btn === none and (select_i !== none)) |=> ##[0:3] select_i !== none)5�_�  '  )          (   �   ,    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      i                       ((inf.flavor_btn === none and (select_i !== none)) |=> (##[0:3] select_i !== none)5�_�  (  +          )   �   ,    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �      m                       ((inf.flavor_btn !== none && inf.flavor_btn !== user_define ) and (select_i === none))5�_�  )  ,  *      +   �   W    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�`     �   �   �   �      n                       ((inf.flavor_btn === no_coffee and (select_i !== none)) |=> (##[0:3] select_i !== none)5�_�  +  -          ,   �   e    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�e     �   �   �   �      n                       ((inf.flavor_btn === no_coffee and (select_i !== none)) |=> (##[1:3] select_i !== none)5�_�  ,  .          -   �       ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4��     �   �   �   �          endproperty5�_�  -  /          .   �        ����                                                                                                                =                                                                                                                                                                                                          �   !       �          V   !    Z4��     �   �   �   �    �   �   �   �    5�_�  .  0          /   �   :    ����                                                                                                                =                                                                                                                                                                                                          �   !       �          V   !    Z4��     �   �   �   �      O    out_valid_cycle_check_general_coffee: assert property(spec5_general_coffee)5�_�  /  1          0   �   1    ����                                                                                                                =                                                                                                                                                                                                          �   1       �   >          >    Z4��     �   �   �   �      �                                $display( "After flavor_btn or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�  0  2          1   �   <    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   U          U    Z4�     �   �   �   �      �                                $display( "After flavor_btn or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�  1  3          2   �   <    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�     �   �   �   �      r                                $display( "After flavor_btn  is high, the out_valid should be high in 30 cycle.");5�_�  2  4          3   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�
     �   �   �   �      j                                $display( "After flavor_btn , the out_valid should be high in 30 cycle.");5�_�  3  5          4   �   =    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�     �   �   �   �      m                                $display( "After flavor_btn () , the out_valid should be high in 30 cycle.");5�_�  4  6          5   �   (    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�     �   �   �   �      G    out_valid_cycle_check_general_coffee: assert property(spec5_supply)5�_�  5  7          6   �        ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�,     �   �   �   �      "                                  �   �   �   �    5�_�  6  8          7   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�;     �   �   �   �              �   �   �   �    5�_�  7  9          8   �   	    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�F     �   �   �   �      	        @5�_�  8  :          9   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�X     �   �   �   �              @(negedge clk)5�_�  9  ;          :   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�X     �   �   �   �              @(negedge clk) 5�_�  :  <          ;   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�X     �   �   �   �              @(negedge clk) ()5�_�  ;  =          <   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�Z     �   �   �   �              @(negedge clk) ()5�_�  <  >          =   �   &    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�]     �   �   �   �      &        @(negedge clk) (inf.out_valid)5�_�  =  ?          >   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�r     �   �   �   �      +        @(negedge clk) (inf.out_valid) ##1 5�_�  >  @          ?   �   ,    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�r     �   �   �   �      -        @(negedge clk) (inf.out_valid) ##1 ()5�_�  ?  A          @   �   ,    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�t     �   �   �   �      -        @(negedge clk) (inf.out_valid) ##1 ()5�_�  @  B          A   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�z     �   �   �   �      ;        @(negedge clk) (inf.out_valid) ##1 (!inf.out_valid)5�_�  A  C          B   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �          �   �   �   �    5�_�  B  D          C   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      I    out_valid_cycle_check_user_define: assert property(spec5_user_define)5�_�  C  E          D   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      ?    out_valid_cycle_check_supply: assert property(spec5_supply)5�_�  D  F          E   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      O    out_valid_cycle_check_general_coffee: assert property(spec5_general_coffee)5�_�  E  G          F   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �          out_valid_1_cycle_check;5�_�  F  H          G   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �          out_valid_1_cycle_check:5�_�  G  I          H   �   #    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      #    out_valid_1_cycle_check: assert5�_�  H  J          I   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      %    out_valid_1_cycle_check: assert()5�_�  I  K          J   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      %    out_valid_1_cycle_check: assert()5�_�  J  L          K   �   *    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      *    out_valid_1_cycle_check: assert(spec6)5�_�  K  M          L   �   &    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      !                                 �   �   �   �    5�_�  L  N          M   �       ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      !                                 �   �   �   �    5�_�  M  O          N   �   )    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      )                                 $display5�_�  N  P          O   �   *    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      +                                 $display()5�_�  O  Q          P   �   *    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      +                                 $display()5�_�  P  R          Q   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      -                                 $display("")5�_�  Q  S          R   �   ;    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      ;                                 $display("Spec6 is wrong")5�_�  R  T          S   �   )    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      )                                 $display5�_�  S  U          T   �   *    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      +                                 $display()5�_�  T  V          U   �   *    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      +                                 $display()5�_�  U  W          V   �   +    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      -                                 $display("")5�_�  V  X          W   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��    �   �   �   �      "                                  �   �   �   �    5�_�  W  Y          X   �   /    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      <                                 $display("Spec6 is wrong");5�_�  X  Z          Y   �   .    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �      ;                                $display("Spec5 is wrong");5�_�  Y  [          Z   �   .    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�     �   �   �   �      ;                                $display("Spec5 is wrong");5�_�  Z  \          [   �   7    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�     �   �   �   �      D                                         $display("Spec5 is wrong");5�_�  [  ]          \   �   $    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�     �   �   �   �      1                      $display("Spec4 is wrong");5�_�  \  ^          ]   �   2    ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4�    �   �   �   �      ?                                    $display("Spec3 is wrong");5�_�  ]              ^   �        ����                                                                                                                =                                                                                                                                                                                                          �   <       �   C          C    Z4��     �   �   �   �       5�_�  )          +  *   �   W    ����                                                                                                                =                                                                                                                                                                                                          �   4       �   S          S    Z4�P     �   �   �   �      n                       ((inf.flavor_btn === no_coffee and (select_i !== none)) |=> (##[1:3] select_i !== none)5�_�                 �       ����                                                                                                                =                                                                                                                                                                                                          �   @       �   F          F    Z4�&     �   �   �   �          property spec5_;5�_�  
               �   @    ����                                                                                                                =                                                                                                                                                                                                          �   R       �   X          X    Z4�     �   �   �   �      A    out_valid_cycle_check_general_coffee: assert property(spec5_)5�_�                 �   R    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      R                                         $display( "After flavor_btn==user_define 5�_�  �              �   :    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                                         $display( "After (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�                  �   :    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                                         $display( "After also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�                   �   :    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                                         $display( "After depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle.");5�_�  �      �  �  �   �   )    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�L     �   �   �   �    �   �   �   �      "After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle."5�_�  �          �  �   �   (    ����                                                                                                                =                                                                                                                                                                                                          �           �   f              Z4�I     �   �   �   �    �   �   �   �      "After flavor_btn (also depends on ratio signal) or select_i (the last one) is high, the out_valid should be high in 30 cycle."5�_�  i          k  j   �       ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4�0     �   �   �        5�_�            	     �   :    ����                                                                                                                =                                                                                                                                                                                                          �          �                 Z4��     �   �   �   �      �                        if(inf.flavor_out===no_coffee) and(inf.window.espresso.led === red && inf.window.espresso.monitor == 0) and5�_�  �          �  �   �        ����                                                                                                                =                                                                                                                                                                                                          �   ,       �   6          -    Z4�     �   �   �        5�_�  q          s  r   z   
    ����                                                                                                                =                                                                                                                                                                                                          �   .       �   <          <    Z4~�     �   y   {   �      <        @(negedge clk) inf.select_i != 0 |-> inf.supply !=0;5�_�  #          %  $   v        ����                                                                                                                =                                                                                                                                                                                                          v           v           V        Z4wf     �   u   y        5�_�  �  �      �  �   .       ����                                                                                                                <                                                                                                                                                                                                          +          +          V       Z2��     �   -   /        5�_�  �  �          �   .        ����                                                                                                                ;                                                                                                                                                                                                          +          +          V       Z2��     �   -   /        5�_�  �  �          �   .        ����                                                                                                                :                                                                                                                                                                                                          +          +          V       Z2��     �   -   /        5�_�  �              �   .        ����                                                                                                                9                                                                                                                                                                                                          +          +          V       Z2��     �   -   /        5�_�  F          H  G   0       ����                                                                                                                9                                                                                                                                                                                                          ,           .                 Z2�E     �   /   1   f      !    : coverpoint inf.flavor_btn{ 5�_�   �              �   K   
    ����                                                                                                                7                                                                                                                                                                                                          G          G   #          #    Z2��     �   J   M   ]      ,        bins inf.window.milk.led{ = {green};5�_�   �           �   �   N       ����                                                                                                                7                                                                                                                                                                                                          F          Q                 Z2�s     �   N   O   X       5�_�   �       �   �   �   F       ����                                                                                                                7                                                                                                                                                                                                          F          J                 Z2��     �   F   G   N    �   F   G   N          option.per_instance = 1;5�_�   �           �   �   F       ����                                                                                                                7                                                                                                                                                                                                          F          I                 Z2��     �   E   G   N      3    bins espresso_led  : {inf.window.espresso.led};�   F   J   N      /    bins milk_led      : {inf.window.milk.led};   4    bins chocolate_led : {inf.window.chocolate.led};   0    bins froth_led     : {inf.window.froth.led};5��