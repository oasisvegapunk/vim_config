Vim�UnDo� �gr����L����#Ӳ�K;9�R� �`��y   (                 ^       ^   ^   ^    Z��    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Z�{     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʂ     �                  module FP_add5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʂ     �                  module FP_add()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʃ     �                  module FP_add()5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             Zʏ    �                  *module FP_add(ae, am, be, bm, ce, cm, ovf)5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             Zʑ    �                  �               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʗ     �               �               5�_�      	                 
    ����                                                                                                                                                                                                                                                                                                                                                             Zʚ     �                 parameter e =3;5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             Zʜ     �                 parameter m =3;5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             Zʝ     �                  �               5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             Zʟ     �                �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʤ     �               input 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʨ     �               input [e-1:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʨ    �               input [e-1:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʭ     �             �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             Zʭ     �             �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʲ     �               input [e-1:0] ae, be;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             Zʶ     �               input [e-1:0] ae, be;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʸ     �               output[e-1:0] ae, be;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʺ     �      	   	       �      	       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Zʼ     �      	   	      output 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �      	   	      output [m-1:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��    �      	   	      output [m-1:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �      	   	      output [m-1:0] am,bm;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �      	   	      output [m-1:0] ;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         	      output [e-1:0] ae, be;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��    �         	      output [e-1:0] ;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         	      input [e-1:0] ae, be;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         	      input [m-1:0] ae, be;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         	      output [e-1:0] ce;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             Z��    �      	   	      output [m-1:0] cm;5�_�      !                  $    ����                                                                                                                                                                                                                                                                                                                                                             Z̟     �      
   
       �      
   	    5�_�       "           !   	        ����                                                                                                                                                                                                                                                                                                                                                             Z̬     �   	             �   	      
    5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                             Z̰     �   
             5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             Z̲     �   
            wire 5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                             Z̲     �   
            wire []5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             Z̳     �   
            wire []5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             Z̶    �   
            wire [e-1:0]5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                             Z̽     �                �             5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             Z̿     �               wire 5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             Z̿     �               wire []5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               wire []5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             Z��    �               wire [m-1:0]5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             Z��   	 �                �             5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                �             5�_�   -   /           .           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               wire agtb = 5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               wire agtb = ()5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               wire agtb = ()5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               wire agtb = (ae >= be)5�_�   2   4           3      *    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                �             5�_�   3   5           4      .    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �             �             5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               /assign ge = agtb ? ae : be; // greater exponent5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                             Z�      �               /assignlge = agtb ? ae : be; // greater exponent5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �               /assign le = agtb ? ae : be; // greater exponent5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �               /assign le = agtb ? be : be; // greater exponent5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                             Z�   
 �               /assign le = agtb ? be : ae; // greater exponent5�_�   9   ;           :      &    ����                                                                                                                                                                                                                                                                                                                                                             Z�    �                �             5�_�   :   <           ;      *    ����                                                                                                                                                                                                                                                                                                                                                             Z�,    �                �             5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                             Z�G     �                �             5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                             Z�T     �               assign gm = agtb ? am : bm;5�_�   =   ?           >      #    ����                                                                                                                                                                                                                                                                                                                                                             Z�Z    �               /assign gm = agtb ? am : bm; // greter mantissas5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                             Z�a    �               assign lm = agtb ? bm : am; 5�_�   ?   A           @      /    ����                                                                                                                                                                                                                                                                                                                                                             Z�i     �                �             5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                             Z�o     �               // �             5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                             Z͈    �               assign alm = lm >> de;5�_�   B   D           C      9    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               9assign alm = lm >> de;// align mantissas with smaller one5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               )assign alm = lm >> de;// align mantissas 5�_�   D   F           E      1    ����                                                                                                                                                                                                                                                                                                                                                             Z��    �               1assign alm = lm >> de;// align smaller mantissas 5�_�   E   G           F      >    ����                                                                                                                                                                                                                                                                                                                                                             Z��    �                �             5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                // find first one5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                             Z�
    �         !      sc // shift cound5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �      !   "       �          !    5�_�   I   K           J           ����                                                                                                                                                                                                                                                                                                                                                             Z�     �      !   #      assign 5�_�   J   L           K           ����                                                                                                                                                                                                                                                                                                                                                             Z�     �      !   #      	assign {}5�_�   K   M           L           ����                                                                                                                                                                                                                                                                                                                                                             Z�     �      !   #      	assign {}5�_�   L   N           M           ����                                                                                                                                                                                                                                                                                                                                                             Z�     �      !   #      assign {nm,rnd}5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                                                             Z�)     �         $       �         #    5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                                                             Z�,     �         %      wire 5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                                                             Z�,     �         %      wire []5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                                             Z�-     �         %      wire []5�_�   Q   S           R      
    ����                                                                                                                                                                                                                                                                                                                                                             Z�0    �         %      
wire [m:0]5�_�   R   T           S           ����                                                                                                                                                                                                                                                                                                                                                             Z�E     �      !   %      sc // shift count5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                             Z�H    �          %      // find first one5�_�   T   V           U   "       ����                                                                                                                                                                                                                                                                                                                                                             Z�[    �   !   #   %      assign {nm,rnd} = sm << 5�_�   U   W           V   "       ����                                                                                                                                                                                                                                                                                                                                                             Z�^     �   "   $   &       �   "   $   %    5�_�   V   X           W   #       ����                                                                                                                                                                                                                                                                                                                                                             Z�`     �   "   $   &      assign 5�_�   W   Y           X   #       ����                                                                                                                                                                                                                                                                                                                                                             Z�`     �   "   $   &      	assign {}5�_�   X   Z           Y   #       ����                                                                                                                                                                                                                                                                                                                                                             Z�a     �   "   $   &      	assign {}5�_�   Y   [           Z   #       ����                                                                                                                                                                                                                                                                                                                                                             Z�c    �   "   $   &      assign {ovf,ce}5�_�   Z   \           [   #   7    ����                                                                                                                                                                                                                                                                                                                                                             Z��    �   #   &   '       �   #   %   &    5�_�   [   ]           \   %       ����                                                                                                                                                                                                                                                                                                                                                             Z��    �   %   '   )      // �   %   '   (    5�_�   \   ^           ]   &        ����                                                                                                                                                                                                                                                                                                                                                             Z��    �   %   '   )      // assign cm = nm + rnd;5�_�   ]               ^   '        ����                                                                                                                                                                                                                                                                                                                                                             Z��    �   &   '           5��