Vim�UnDo� �r���8��y?`��6��|ۈ�*�|�P  q              �  �      �  �  �    Z"X�   M _�       �           �   Y       ����                                                                                                                                                                                                                                                                                                                            X          \                 Z �"     �   X   Z   b      .            S_GENERAL_REQ: espresso_weight <= 5�_�   �   �           �   Y       ����                                                                                                                                                                                                                                                                                                                            X          \                 Z �#     �   X   [   b      .            S_GENERAL_REQ: espresso_weight <= 5�_�   �   �           �   Y       ����                                                                                                                                                                                                                                                                                                                            X          ]                 Z �%     �   Y   [   d                      �   Y   [   c    5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            X          ^                 Z �'     �   Y   [   d                      case5�_�   �   �           �   Z   "    ����                                                                                                                                                                                                                                                                                                                            X          ^                 Z �/     �   Y   [   d      #                case(required_size)5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            X          ^                 Z �2     �   [   ]   e                          �   [   ]   d    5�_�   �   �   �       �   Z       ����                                                                                                                                                                                                                                                                                                                            X          _                 Z �;     �   Y   [   e      #                case(required_size)5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            X          _                 Z �R     �   Z   \   e      #                espresso_weight <= 5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            X          _                 Z �S     �   Z   \   e      #                espresso_weight <= 5�_�   �              �   [       ����                                                                                                                                                                                                                                                                                                                            X          _                 Z �V     �   Z   \   e      '                    espresso_weight <= 5�_�   �                [       ����                                                                                                                                                                                                                                                                                                                            X          _                 Z �X     �   Z   \   e      (                    :espresso_weight <= 5�_�                  [       ����                                                                                                                                                                                                                                                                                                                            X          _                 Z �Z     �   [   ]   f                              �   [   ]   e    5�_�                 U       ����                                                                                                                                                                                                                                                                                                                            X          `                 Z �i     �   U   W   g              �   U   W   f    5�_�                 V       ����                                                                                                                                                                                                                                                                                                                            Y          a                 Z �o     �   U   W   g              milk_weight <= 5�_�                 V       ����                                                                                                                                                                                                                                                                                                                            Y          a                 Z �p     �   U   W   g              milk_weight <= 'b0'5�_�                 V       ����                                                                                                                                                                                                                                                                                                                            Y          a                 Z �q     �   U   W   g              milk_weight <= 'b0'5�_�                 V       ����                                                                                                                                                                                                                                                                                                                            Y          a                 Z �r     �   V   X   h              �   V   X   g    5�_�                 W       ����                                                                                                                                                                                                                                                                                                                            Z          b                 Z �{     �   V   X   h              chocolate_weight <= 5�_�    	             W       ����                                                                                                                                                                                                                                                                                                                            Z          b                 Z �|     �   V   X   h               chocolate_weight <= 'b0'5�_�    
          	   W        ����                                                                                                                                                                                                                                                                                                                            Z          b                 Z �}     �   V   X   h               chocolate_weight <= 'b0'5�_�  	            
   W       ����                                                                                                                                                                                                                                                                                                                            Z          b                 Z �~     �   W   Y   i              �   W   Y   h    5�_�  
               X       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z Ë     �   W   Y   i              froth_weight  <= 5�_�                 X       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z Ì     �   W   Y   i              froth_weight  <= 'b0'5�_�                 X       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z Ì     �   W   Y   i              froth_weight  <= 'b0'5�_�                 X       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z Ð     �   W   Y   i              froth_weight  <= 'b0;5�_�                 V       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z Ó     �   U   W   i              milk_weight <= 'b0;5�_�                 U       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z Ö     �   T   V   i              espresso_weight <= 'b0;5�_�                 ^       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z Þ     �   ]   _   i      -                    latte:espresso_weight <= 5�_�                 ^       ����                                                                                                                                                                                                                                                                                                                            [          c                 Z ß     �   ]   _   i      -                    latte:espresso_weight <= 5�_�                 ^        ����                                                                                                                                                                                                                                                                                                                            [          c                 Z á     �   ]   `   i      3                    latte: beginespresso_weight <= 5�_�                 _   +    ����                                                                                                                                                                                                                                                                                                                            [          d                 Z ��     �   ^   `   j      +                        espresso_weight <= 5�_�                 _   ,    ����                                                                                                                                                                                                                                                                                                                            [          d                 Z ��     �   ^   `   j      ,                        espresso_weight <= 45�_�                 _        ����                                                                                                                                                                                                                                                                                                                            U          X           V   /    Z ��     �   _   d   j    �   _   `   j    5�_�                 `       ����                                                                                                                                                                                                                                                                                                                            `          c                 Z ��     �   `   d   n               milk_weight      <= 'b0;            chocolate_weight <= 'b0;            froth_weight     <= 'b0;�   _   a   n               espresso_weight  <= 'b0;5�_�                 `   
    ����                                                                                                                                                                                                                                                                                                                            `          c                 Z ��     �   _   `          0                        espresso_weight  <= 'b0;5�_�                 `   -    ����                                                                                                                                                                                                                                                                                                                            `   -       b   -          -    Z ��     �   _   c   m      0                        milk_weight      <= 'b0;   0                        chocolate_weight <= 'b0;   0                        froth_weight     <= 'b0;5�_�                 `   +    ����                                                                                                                                                                                                                                                                                                                            `   +       b   +          +    Z ��     �   _   c   m      0                        milk_weight      <= 'd0;   0                        chocolate_weight <= 'd0;   0                        froth_weight     <= 'd0;5�_�                 `   .    ����                                                                                                                                                                                                                                                                                                                            `   +       b   +          +    Z ��     �   _   a   m      0                        milk_weight      <=4'd0;5�_�                 b   .    ����                                                                                                                                                                                                                                                                                                                            `   +       b   +          +    Z ��     �   a   c   m      0                        froth_weight     <=4'd0;5�_�                 b   .    ����                                                                                                                                                                                                                                                                                                                            `   +       b   +          +    Z ��     �   b   d   n                              �   b   d   m    5�_�                 c       ����                                                                                                                                                                                                                                                                                                                            `   +       b   +          +    Z ��     �   c   e   o                          �   c   e   n    5�_�                  d   #    ����                                                                                                                                                                                                                                                                                                                            `   +       b   +          +    Z ��     �   d   f   p                              �   d   f   o    5�_�    !              d       ����                                                                                                                                                                                                                                                                                                                            `   +       b   +          +    Z ��     �   d   f   p    5�_�     "          !   d        ����                                                                                                                                                                                                                                                                                                                            _          b          V       Z ��     �   d   i   q    �   d   e   q    5�_�  !  #          "   i        ����                                                                                                                                                                                                                                                                                                                            _          b          V       Z ��     �   h   i           5�_�  "  $          #   h   .    ����                                                                                                                                                                                                                                                                                                                            _          b          V       Z ��     �   g   i   t      0                        froth_weight     <=4'd2;5�_�  #  %          $   i       ����                                                                                                                                                                                                                                                                                                                            _          b          V       Z �     �   i   k   u                          �   i   k   t    5�_�  $  &          %   j       ����                                                                                                                                                                                                                                                                                                                            _          b          V       Z �     �   j   l   v                              �   j   l   u    5�_�  %  '          &   j       ����                                                                                                                                                                                                                                                                                                                            _          b          V       Z �     �   j   l   v    �   j   k   v    5�_�  &  (          '   j        ����                                                                                                                                                                                                                                                                                                                            e           h           V        Z �     �   j   o   w    �   j   k   w    5�_�  '  )          (   o        ����                                                                                                                                                                                                                                                                                                                            e           h           V        Z �     �   n   o           5�_�  (  *          )   _   +    ����                                                                                                                                                                                                                                                                                                                            _   +       b   +          +    Z �'     �   ^   c   z      0                        espresso_weight <= 4'd2;   0                        milk_weight      <=4'd1;   0                        chocolate_weight <=4'd0;   0                        froth_weight     <=4'd2;5�_�  )  +          *   e   +    ����                                                                                                                                                                                                                                                                                                                            e   +       h   +          +    Z �)     �   d   i   z      0                        espresso_weight <= 4'd2;   0                        milk_weight      <=4'd1;   0                        chocolate_weight <=4'd0;   0                        froth_weight     <=4'd1;5�_�  *  ,          +   k   +    ����                                                                                                                                                                                                                                                                                                                            k   +       n   +          +    Z �-     �   j   o   z      0                        espresso_weight <= 4'd2;   0                        milk_weight      <=4'd1;   0                        chocolate_weight <=4'd0;   0                        froth_weight     <=4'd1;5�_�  +  -          ,   k   .    ����                                                                                                                                                                                                                                                                                                                            k   +       n   +          +    Z �3     �   j   l   z      0                        espresso_weight <= 3'd2;5�_�  ,  .          -   m   .    ����                                                                                                                                                                                                                                                                                                                            k   +       n   +          +    Z �4     �   l   n   z      0                        chocolate_weight <=3'd0;5�_�  -  /          .   n   .    ����                                                                                                                                                                                                                                                                                                                            k   +       n   +          +    Z �5     �   m   o   z      0                        froth_weight     <=3'd1;5�_�  .  0          /   R       ����                                                                                                                                                                                                                                                                                                                            k   +       n   +          +    Z �?     �   Q   S   z      logic [3:0] espresso_weight;5�_�  /  1          0   R       ����                                                                                                                                                                                                                                                                                                                            k   +       n   +          +    Z �A     �   R   T   z    �   R   S   z    5�_�  0  2          1   R       ����                                                                                                                                                                                                                                                                                                                            V          Y                 Z �I     �   R   T   {    5�_�  1  3          2   T        ����                                                                                                                                                                                                                                                                                                                            W          Z                 Z �K     �   S   X   |       5�_�  2  4          3   S        ����                                                                                                                                                                                                                                                                                                                            Z          ]                 Z �M     �   R   X                          �   S   T       5�_�  3  5          4   R       ����                                                                                                                                                                                                                                                                                                                            Z          ]                 Z �T     �   Q   S         logic [2:0] espresso_weight;5�_�  4  6          5   R       ����                                                                                                                                                                                                                                                                                                                            Z          ]                 Z �U     �   Q   S         logic [2:0]    espresso_weight  5�_�  5  7          6   R       ����                                                                                                                                                                                                                                                                                                                            Y          \                 Z �W     �   Q   S   ~      logic [2:0] espresso_weight  5�_�  6  8          7   S       ����                                                                                                                                                                                                                                                                                                                            Y          \                 Z �\     �   R   T   ~      milk_weight      5�_�  7  9          8   T       ����                                                                                                                                                                                                                                                                                                                            Y          \                 Z �_     �   S   U   ~      chocolate_weight 5�_�  8  :          9   U       ����                                                                                                                                                                                                                                                                                                                            Y          \                 Z �a     �   T   V   ~      froth_weight     5�_�  9  ;          :   S        ����                                                                                                                                                                                                                                                                                                                            S           U                   Z �g     �   S   V   ~      chocolate_weight,   froth_weight;�   R   T   ~      milk_weight,     5�_�  :  <          ;   s        ����                                                                                                                                                                                                                                                                                                                            S           U                   Z ă     �   s   u                             �   s   u   ~    5�_�  ;  =          <   t        ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z Ĕ     �   t   y       �   t   u       5�_�  <  >          =   u   .    ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ė     �   t   v   �      0                        espresso_weight <= 3'd1;5�_�  =  ?          >   v   .    ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ę     �   u   w   �      0                        milk_weight      <=3'd1;5�_�  >  @          ?   w   .    ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z Ě     �   v   x   �      0                        chocolate_weight <=3'd1;5�_�  ?  A          @   x   .    ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ě     �   w   y   �      0                        froth_weight     <=3'd0;5�_�  @  B          A   y        ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ��     �   x   y           5�_�  A  C          B   {       ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ��     �   z   {          0            S_CUSTOMIZED_REQ: espresso_weight <=5�_�  B  D          C   y       ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ��     �   y   |   �                      �   y   {   �    5�_�  C  E          D   z       ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ��     �   y   {   �                  S_MILK:5�_�  D  F          E   {       ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z ��     �   {   ~   �                  �   {   }   �    5�_�  E  G          F   z       ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z �)     �   y   {   �                  S_ESPRESSO:5�_�  F  H          G   z       ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z �+     �   z   |   �                          �   z   |   �    5�_�  G  I          H   z       ����                                                                                                                                                                                                                                                                                                                            o          r          V       Z �-     �   z   |   �    5�_�  H  J          I   z        ����                                                                                                                                                                                                                                                                                                                            u          x          V       Z �3     �   z      �    �   z   {   �    5�_�  I  K          J           ����                                                                                                                                                                                                                                                                                                                            u          x          V       Z �5     �   ~              5�_�  J  L          K   {   /    ����                                                                                                                                                                                                                                                                                                                            u          x          V       Z �9     �   z   |   �      0                        espresso_weight <= 3'd0;5�_�  K  M          L   {   (    ����                                                                                                                                                                                                                                                                                                                            u          x          V       Z �A     �   z   |   �      1                        espresso_weight <= ratio;5�_�  L  N          M   |   +    ����                                                                                                                                                                                                                                                                                                                            |   +       ~   .          .    Z �E     �   {      �      0                        milk_weight      <=3'd0;   0                        chocolate_weight <=3'd0;   0                        froth_weight     <=3'd0;5�_�  M  O          N   |   *    ����                                                                                                                                                                                                                                                                                                                            |          ~   (          (    Z �N     �   {   �   �      ,                        milk_weight      <=;   ,                        chocolate_weight <=;   ,                        froth_weight     <=;                   end�   |   }   �    5�_�  N  P          O   |   +    ����                                                                                                                                                                                                                                                                                                                            |   +       ~   +          +    Z �P     �   |      �      =                        chocolate_weight <=chocolate_weight ;   =                        froth_weight     <=froth_weight     ;�   {   }   �      =                        milk_weight      <=milk_weight      ;5�_�  O  Q          P   |   <    ����                                                                                                                                                                                                                                                                                                                            |   <       ~   <          <    Z �T     �   {      �      >                        milk_weight      <= milk_weight      ;   >                        chocolate_weight <= chocolate_weight ;   >                        froth_weight     <= froth_weight     ;5�_�  P  R          Q   �       ����                                                                                                                                                                                                                                                                                                                            |   <       ~   <          <    Z �X     �      �   �                  S_MILK:5�_�  Q  S          R   �       ����                                                                                                                                                                                                                                                                                                                            |   <       ~   <          <    Z �Y     �   �   �   �                          �   �   �   �    5�_�  R  T          S   z       ����                                                                                                                                                                                                                                                                                                                            |   <       ~   <          <    Z �q     �   y   {   �                       S_ESPRESSO:begin5�_�  S  U          T   �       ����                                                                                                                                                                                                                                                                                                                            |   <       ~   <          <    Z �s     �      �   �                      S_MILK:begin5�_�  T  V          U   �        ����                                                                                                                                                                                                                                                                                                                            u          x          V       Z ŀ     �   �   �   �    �   �   �   �    5�_�  U  W          V   �   (    ����                                                                                                                                                                                                                                                                                                                            u          x          V       Z ń     �   �   �   �      0                        espresso_weight <= 3'd0;5�_�  V  X          W   �   +    ����                                                                                                                                                                                                                                                                                                                            �   +       �   +          +    Z Ŋ     �   �   �   �      0                        chocolate_weight <=3'd0;   0                        froth_weight     <=3'd0;�   �   �   �      0                        milk_weight      <=3'd0;5�_�  W  Y          X   �   ,    ����                                                                                                                                                                                                                                                                                                                            �   ,       �   /          /    Z ō     �   �   �   �      1                        espresso_weight  <= 3'd0;   1                        milk_weight      <= 3'd0;   1                        chocolate_weight <= 3'd0;   1                        froth_weight     <= 3'd0;5�_�  X  Z          Y   �   +    ����                                                                                                                                                                                                                                                                                                                            �          �   '          '    Z Ŕ     �   �   �   �      -                        espresso_weight  <= ;   -                        milk_weight      <= ;   -                        chocolate_weight <= ;   -                        froth_weight     <= ;                   end�   �   �   �    5�_�  Y  [          Z   �        ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z ś     �   �   �   �    �   �   �   �    5�_�  Z  \          [   �       ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z Ŝ     �   �   �   �                  S_CHOCOLATE:5�_�  [  ]          \   �        ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z ş     �   �   �   �                              �   �   �   �    5�_�  \  ^          ]   �       ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z ţ     �   �   �   �      !                S_CHOCOLATE:begin5�_�  ]  _          ^   �       ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z Ŧ     �   �   �   �                          end5�_�  ^  `          _   �       ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z Ũ     �   �   �   �                  S_FROTH:5�_�  _  a          `   �       ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z Ū     �   �   �   �                          �   �   �   �    5�_�  `  c          a   �       ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z ŭ     �   �   �   �                      S_FROTH:begin5�_�  a  d  b      c   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ŵ     �   �   �   �    �   �   �   �    5�_�  c  e          d   �   ,    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ź     �   �   �   �      =                        milk_weight      <= milk_weight     ;5�_�  d  f          e   {   ,    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   z   |   �      2                        espresso_weight  <= ratio;5�_�  e  g          f   �   ,    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �      2                        milk_weight      <= ratio;5�_�  f  h          g   �   +    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �      =                        chocolate_weight <= chocolate_weight;5�_�  g  i          h   �   ,    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �      =                        froth_weight     <= froth_weight    ;5�_�  h  j          i   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �      6                        froth_weight     <= inf.ratio;5�_�  i  k          j   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �      =                        froth_weight     <= inf.ratio       ;5�_�  j  l          k   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �                      �   �   �   �    5�_�  k  m          l   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �                  default:�   �   �   �    5�_�  l  n          m   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �                  default:       5�_�  m  o          n   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �                      �   �   �   �    5�_�  n  p          o   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �     �   �   �   �      #                default:begin      5�_�  o  q          p   `       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �     �   _   a   �                  S_GENERAL_REQ: 5�_�  p  r          q   y       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �     �   y   {   �                      �   y   {   �    5�_�  q  s          r   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �     �   �   �   �    �   �   �   �    5�_�  r  t          s   �   ,    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �     �   �   �   �      6                        froth_weight     <= inf.ratio;5�_�  s  u          t   �   ,    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �     �   �   �   �      -                        froth_weight     <= ;5�_�  t  v          u   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �/     �   �   �           5�_�  u  w          v   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �Y     �   �   �   �       �   �   �   �    5�_�  v  x          w   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �]     �   �   �   �      logic 5�_�  w  y          x   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �]     �   �   �   �      logic []5�_�  x  z          y   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �t     �   �   �   �      logic []5�_�  y  {          z   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �y     �   �   �   �      logic [4:0]5�_�  z  |          {   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƀ     �   �   �   �       �   �   �   �    5�_�  {  }          |   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ƈ     �   �   �   �      assign sum_weight = 5�_�  |  ~          }   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƈ     �   �   �   �      assign sum_weight = ()5�_�  }            ~   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ɖ     �   �   �   �      assign sum_weight = ()5�_�  ~  �             �   8    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ǝ     �   �   �   �      8assign sum_weight = (espresso_weight + chocolate_weight)5�_�    �          �   �   ;    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ɛ     �   �   �   �      ;assign sum_weight = (espresso_weight + chocolate_weight) + 5�_�  �  �          �   �   <    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ɛ     �   �   �   �      =assign sum_weight = (espresso_weight + chocolate_weight) + ()5�_�  �  �          �   �   &    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ɩ     �   �   �   �      =assign sum_weight = (espresso_weight + chocolate_weight) + ()5�_�  �  �          �   �   7    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƚ     �   �   �   �      8assign sum_weight = (espresso_weight + milk_weight) + ()5�_�  �  �          �   �   W    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ơ   	 �   �   �   �      Wassign sum_weight = (espresso_weight + milk_weight) + (chocolate_weight + froth_weight)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƣ     �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ƥ     �   �   �           5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƥ     �   �   �   �       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƴ     �   �   �   �      logic 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƴ     �   �   �   �      logic []5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ƽ     �   �   �   �      logic []5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �      logic [] user_define_basis;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �      logic [9:0] user_define_basis;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z ��     �   �   �   �       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �   
 �   �   �   �      assign user_define_basis = 5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �4     �   �   �          logic [9:0] user_define_basis;5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �5     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �7     �   �   �          logic [9:0] user_define_basis;5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �8     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �;     �   �   �   �       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �C     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �D     �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �e     �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �$    �   �   �   �       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �W     �   �   �   �      /// This should change to the accumulate version5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �Z     �   �   �   �       �   �   �   �    5�_�  �  �          �   �   3    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �_     �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �`     �   �   �          //5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �a     �   �   �   �      //�   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �k     �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �n     �   �   �   �       �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z Ȫ     �   �   �   �       5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            M          P          V       Z ��     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      logic [9:0] espresso_req;   logic [9:0] milk_req;   logic [9:0] chocolate_req;   logic [9:0] froth_req;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      espresso_req;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      	milk_req;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      chocolate_req;5�_�  �  �          �   �   	    ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      
froth_req;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      espresso_req5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      espresso_req = ingredient_basis5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      begin5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �     �   �   �   �      begin if5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �     �   �   �   �      espresso_req = ingredient_basis5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �     �   �   �   �      milk_req5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �"     �   �   �   �       milk_req     = ingredient_base *5�_�  �  �          �   �   !    ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �#     �   �   �   �      !milk_req     = ingredient_base  *5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �(     �   �   �   �      chocolate_req5�_�  �  �          �   �   	    ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �0     �   �   �   �      	froth_req5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �4     �   �   �   �      froth_req   = 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �5     �   �   �   �      froth_req    = 5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �>     �   �   �           5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �C     �   �   �   �      2espresso_req = ingredient_basis * espresso_weight;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �D     �   �   �   �      .milk_req     = ingredient_base  * milk_weight;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �E     �   �   �   �      3chocolate_req = ingredient_base * chocolate_weight;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �F     �   �   �   �      0froth_req    = ingredient_base  * froth_weight; 5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �T     �   �   �   �       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �W     �   �   �   �      logic 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �W     �   �   �   �      logic []5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �i     �   �   �   �      logic []5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �m     �   �   �   �      logic [9:0]5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ɉ     �   �   �   �      logic []  ingredient_base = 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ɉ    �   �   �   �      logic []  ingredient_base = ()5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ɪ     �   �   �   �      Elogic []  ingredient_base = () ? user_define_basis : ingredient_base;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ɲ     �   �   �   �      logic [9:0] user_define_basis;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ɳ     �   �   �   �      logic [9:0] user_define_bass;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ɴ     �   �   �   �      logic [9:0] user_define_bas;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ɷ     �   �   �   �      8assign user_define_basis = ingredient_base / sum_weight;5�_�  �  �          �   �   2    ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      Glogic []  ingredient_basis  = () ? user_define_basis : ingredient_base;5�_�  �  �          �   �   2    ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      Flogic []  ingredient_basis  = () ? user_define_bass : ingredient_base;5�_�  �  �          �   �   2    ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      Elogic []  ingredient_basis  = () ? user_define_bas : ingredient_base;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �      Flogic []  ingredient_basis  = () ? user_define_base : ingredient_base;5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��    �   �   �   �      3chocolate_req = ingredient_base * chocolate_weight;5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                 Z ��     �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      4chocolate_req = ingredient_base  * chocolate_weight;   1froth_req     = ingredient_base  * froth_weight; �   �   �   �      /milk_req      = ingredient_base  * milk_weight;5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �      1milk_req      = ingredient_basise  * milk_weight;   6chocolate_req = ingredient_basise  * chocolate_weight;   3froth_req     = ingredient_basise  * froth_weight; 5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �    �   �   �   �      0milk_req      = ingredient_basis  * milk_weight;   5chocolate_req = ingredient_basis  * chocolate_weight;   2froth_req     = ingredient_basis  * froth_weight; 5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �    �   �   �   �       �   �   �   �    5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                                                             Z ̩     �   1   3   �                  weight_size<= 'd0;5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                                                             Z ̪     �   1   3   �                  weight_size <= 'd0;5�_�  �  �          �   ?   	    ����                                                                                                                                                                                                                                                                                                                                                             Z ̰     �   >   @   �          else begin 5�_�  �  �          �   ?       ����                                                                                                                                                                                                                                                                                                                                                             Z ̱     �   >   @   �          else ifbegin 5�_�  �  �          �   ?       ����                                                                                                                                                                                                                                                                                                                                                             Z ̵     �   >   @   �          else if()begin 5�_�  �  �          �   ?       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   >   @   �      #    else if(c_state == INPUT)begin 5�_�  �  �          �   ?       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   >   @   �      %    else if(c_state == S_INPUT)begin 5�_�  �  �          �   A       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   A   C   �          �   A   C   �    5�_�  �  �          �   B       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   B   D   �              �   B   D   �    5�_�  �  �          �   B       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   B   D   �              �   B   D   �    5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   E   G   �    5�_�  �  �          �   L       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   K   M   �          else begin 5�_�  �  �          �   L       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   K   M   �          else if begin 5�_�  �  �          �   L       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   K   M   �      &    else if(n_state == S_INPUT) begin 5�_�  �  �          �   N       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   N   P   �          �   N   P   �    5�_�  �  �          �   O       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   O   Q   �              �   O   Q   �    5�_�  �  �          �   O       ����                                                                                                                                                                                                                                                                                                                                                             Z �      �   O   Q   �              �   O   Q   �    5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   R   T   �    5�_�  �  �          �   :        ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   9   ;   �       5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   R   T   �       �   R   T   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z Ϳ     �   �   �   �       �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   �   �   �       �   �   �   �    5�_�  �  �          �   �   <    ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   �   �   �       �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   �   �   �      //�   �   �   �    5�_�  �  �          �   �   =    ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   �   �   �      =// ---------------- ingredient_basis should be stored -------5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   �   �   �       �   �   �   �    5�_�  �  �          �   �   <    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      //�   �   �   �    5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      =//------------------- COMPARE & UPDATE ----------------------5�_�  �  �          �   �   1    ����                                                                                                                                                                                                                                                                                                                                                             Z �    �   �   �   �      =//-----------------------------------------------------------5�_�  �  �          �   )        ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   )   +   �    5�_�  �  �          �   *        ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �   )   *           5�_�  �  �          �   +       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   *   ,   �      begin: base_selector5�_�  �  �          �   ;   1    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   :   <   �      1always_ff@(posedge clk or negedge inf.rst_n)begin5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z �o     �   �   �           5�_�  �  �          �   �   "    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      Ilogic [9:0]  ingredient_basis  = () ? user_define_base : ingredient_base;5�_�  �  �          �   �   <    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      //�   �   �   �    5�_�  �  �          �   �   
    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      
always_ff@5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      (always_ff@(posedge clk or negedge rst_n)5�_�  �  �          �   �   (    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      (always_ff@(posedge clk or negedge rst_n)5�_�  �  �          �   �   ,    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �          if5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �          if(!inf.rst_n)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �          if(!inf.rst_n)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �              �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �              �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �    5�_�  �             �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �       �   �   �   �    5�_�  �                �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      logic 5�_�                  �   
    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      logic [9:0]5�_�                 �       ����                                                                                                                                                                                                                                                                                                                                                             Z �     �   �   �   �      logic [9:0]5�_�               �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �'     �   �   �   �       �   �   �   �    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �,     �   �   �   �      logic [9:0]                 �   �   �   �    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �/     �   �   �   �      logic [9:0] espresso_req 5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �6     �   �   �   �                  milk_req     5�_�    	             �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �8     �   �   �   �                  milk_rea     5�_�    
          	   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �:     �   �   �   �                  chocolate_req5�_�  	            
   �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �?     �   �   �   �                  froth_req    5�_�  
               �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �E     �   �   �   �      logic [9:0] espresso_remain 5�_�               �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �L     �   �   �   �                  milk_remain     5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �R     �   �   �   �                  chocolate_remain5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z �Z     �   �   �   �    �   �   �   �    5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �_     �   �   �   �      logic [9:0] espresso_remain,5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �b     �   �   �   �                  espresso_remain,5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �c     �   �   �   �                  milk_remain,    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �e     �   �   �   �                  milk_remain, 5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �g     �   �   �   �                  chocolate_remain,5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �i     �   �   �   �                  froth_remain;    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �j     �   �   �   �                  espresso_remain5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �m     �   �   �   �                  espresso_remain5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �r     �   �   �   �                  espresso_remain  5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �s     �   �   �   �                   espresso_remain <=  5�_�                 �   "    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �u     �   �   �   �      $            espresso_remain <= 'b0' 5�_�                 �   $    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �u     �   �   �   �                  milk_remain                chocolate_remain               froth_remain    �   �   �   �      $            espresso_remain <= 'b0' 5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �x     �   �   �           5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �{     �   �   �   �                  milk_remain 5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �                  milk_remain     <= 5�_�                  �   "    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      #            milk_remain     <= 'b0'5�_�    !              �   #    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      #            milk_remain     <= 'b0'5�_�     "          !   �   "    ����                                                                                                                                                                                                                                                                                                                            �   !       �   "          "    Z �     �   �   �   �      "            chocolate_remain<= 'b05�_�  !  #          "   �        ����                                                                                                                                                                                                                                                                                                                            �   "       �   "       V   "    Z �     �   �   �   �    �   �   �   �    5�_�  "  $          #   �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   "       V   "    Z �     �   �   �   �    5�_�  #  %          $   �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   "       V   "    Z �     �   �   �   �              5�_�  $  &          %   �   	    ����                                                                                                                                                                                                                                                                                                                            �   "       �   "       V   "    Z �     �   �   �   �      
        ``5�_�  %  '          &   �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   "       V   "    Z �     �   �   �          
        ``5�_�  &  (          '   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      #            espresso_remain <= 'b0;   #            milk_remain     <= 'b0;   #            chocolate_remain<= 'b0;   "            froth_remain    <= 'b0    �   �   �   �    5�_�  '  )          (   �   /    ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z �     �   �   �   �      3            espresso_remain <= espresso_remain 'b0;   3            milk_remain     <= milk_remain     'b0;   3            chocolate_remain<= chocolate_remain'b0;   2            froth_remain    <= froth_remain    'b05�_�  (  *          )   �   /    ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z �     �   �   �   �      /            froth_remain    <= froth_remain    5�_�  )  +          *   �   "    ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z �     �   �   �   �      "            froth_remain    <= 'b05�_�  *  ,          +   �        ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �           5�_�  +  -          ,   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      0            espresso_remain <= espresso_remain ;5�_�  ,  .          -   �        ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      4            espresso_remain <=(  ) espresso_remain ;5�_�  -  /          .   �   !    ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      5            espresso_remain <=( > ) espresso_remain ;5�_�  .  0          /   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      0            milk_remain     <= milk_remain     ;5�_�  /  1          0   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      2            milk_remain     <=() milk_remain     ;5�_�  0  2          1   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      0            chocolate_remain<= chocolate_remain;5�_�  1  3          2   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      2            chocolate_remain<=() chocolate_remain;5�_�  2  4          3   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �          end5�_�  3  5          4   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      0            froth_remain    <= froth_remain    ;5�_�  4  6          5   �       ����                                                                                                                                                                                                                                                                                                                            �   /       �   1          1    Z ��     �   �   �   �      2            froth_remain    <=() froth_remain    ;5�_�  5  7          6   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      5            espresso_remain <=( > ) espresso_remain ;5�_�  6  8          7   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      4            espresso_remain <=(> ) espresso_remain ;5�_�  7  9          8   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      3            espresso_remain <=( ) espresso_remain ;5�_�  8  :          9   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �	     �   �   �   �      2            espresso_remain <=() espresso_remain ;   2            milk_remain     <=() milk_remain     ;   2            chocolate_remain<=() chocolate_remain;   2            froth_remain    <=() froth_remain    ;           end�   �   �   �    5�_�  9  ;          :   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      B            milk_remain     <=(milk_remain     ) milk_remain     ;   B            chocolate_remain<=(chocolate_remain) chocolate_remain;   B            froth_remain    <=(froth_remain    ) froth_remain    ;�   �   �   �      B            espresso_remain <=(espresso_remain ) espresso_remain ;5�_�  :  <          ;   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      C            espresso_remain <=(>espresso_remain ) espresso_remain ;   C            milk_remain     <=(>milk_remain     ) milk_remain     ;   C            chocolate_remain<=(>chocolate_remain) chocolate_remain;   C            froth_remain    <=(>froth_remain    ) froth_remain    ;5�_�  ;  =          <   �   /    ����                                                                                                                                                                                                                                                                                                                            �   /       �   /          /    Z �      �   �   �   �      B            milk_remain     <=(milk_remain     ) milk_remain     ;   B            chocolate_remain<=(chocolate_remain) chocolate_remain;   B            froth_remain    <=(froth_remain    ) froth_remain    ;�   �   �   �      B            espresso_remain <=(espresso_remain ) espresso_remain ;5�_�  <  >          =   �   /    ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �.     �   �   �   �      D            espresso_remain <=(espresso_remain > ) espresso_remain ;   D            milk_remain     <=(milk_remain     > ) milk_remain     ;   D            chocolate_remain<=(chocolate_remain> ) chocolate_remain;   D            froth_remain    <=(froth_remain    > ) froth_remain    ;           end�   �   �   �    5�_�  =  ?          >   �   0    ����                                                                                                                                                                                                                                                                                                                            �   0       �   0          0    Z �1     �   �   �   �      Q            milk_remain     <=(milk_remain     >milk_req      ) milk_remain     ;   Q            chocolate_remain<=(chocolate_remain>chocolate_req ) chocolate_remain;   Q            froth_remain    <=(froth_remain    >froth_req     ) froth_remain    ;�   �   �   �      Q            espresso_remain <=(espresso_remain >espresso_req  ) espresso_remain ;5�_�  >  @          ?   �   @    ����                                                                                                                                                                                                                                                                                                                            �   @       �   @          @    Z �6     �   �   �   �      R            milk_remain     <=(milk_remain     > milk_req      ) milk_remain     ;   R            chocolate_remain<=(chocolate_remain> chocolate_req ) chocolate_remain;   R            froth_remain    <=(froth_remain    > froth_req     ) froth_remain    ;�   �   �   �      R            espresso_remain <=(espresso_remain > espresso_req  ) espresso_remain ;5�_�  ?  A          @   �       ����                                                                                                                                                                                                                                                                                                                            �   @       �   @          @    Z �F     �   �   �   �              end5�_�  @  B          A   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �W    �   �   �   �      U            milk_remain     <=(milk_remain     > milk_req      )? : milk_remain     ;   U            chocolate_remain<=(chocolate_remain> chocolate_req )? : chocolate_remain;   U            froth_remain    <=(froth_remain    > froth_req     )? : froth_remain    ;�   �   �   �      U            espresso_remain <=(espresso_remain > espresso_req  )? : espresso_remain ;5�_�  A  C          B   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �^    �   �   �           5�_�  B  D          C   �   A    ����                                                                                                                                                                                                                                                                                                                            �           �   >          >    Z �     �   �   �   �      V            espresso_remain <= (espresso_remain > espresso_req  )? : espresso_remain ;   V            milk_remain     <= (milk_remain     > milk_req      )? : milk_remain     ;   V            chocolate_remain<= (chocolate_remain> chocolate_req )? : chocolate_remain;   V            froth_remain    <= (froth_remain    > froth_req     )? : froth_remain    ;       end�   �   �   �    5�_�  C  E          D   �   R    ����                                                                                                                                                                                                                                                                                                                            �   R       �   R          R    Z �     �   �   �   �      u            espresso_remain <= (espresso_remain > espresso_req  )?espresso_remain > espresso_req  : espresso_remain ;   u            milk_remain     <= (milk_remain     > milk_req      )?milk_remain     > milk_req      : milk_remain     ;   u            chocolate_remain<= (chocolate_remain> chocolate_req )?chocolate_remain> chocolate_req : chocolate_remain;   u            froth_remain    <= (froth_remain    > froth_req     )?froth_remain    > froth_req     : froth_remain    ;5�_�  D  F          E   �   B    ����                                                                                                                                                                                                                                                                                                                            �   B       �   B          B    Z �     �   �   �   �      u            milk_remain     <= (milk_remain     > milk_req      )?milk_remain     - milk_req      : milk_remain     ;   u            chocolate_remain<= (chocolate_remain> chocolate_req )?chocolate_remain- chocolate_req : chocolate_remain;   u            froth_remain    <= (froth_remain    > froth_req     )?froth_remain    - froth_req     : froth_remain    ;�   �   �   �      u            espresso_remain <= (espresso_remain > espresso_req  )?espresso_remain - espresso_req  : espresso_remain ;5�_�  E  G          F   �        ����                                                                                                                                                                                                                                                                                                                            �           �   >          >    Z �     �   �   �   �      v            espresso_remain <= (espresso_remain > espresso_req  )? espresso_remain - espresso_req  : espresso_remain ;   v            milk_remain     <= (milk_remain     > milk_req      )? milk_remain     - milk_req      : milk_remain     ;   v            chocolate_remain<= (chocolate_remain> chocolate_req )? chocolate_remain- chocolate_req : chocolate_remain;   v            froth_remain    <= (froth_remain    > froth_req     )? froth_remain    - froth_req     : froth_remain    ;5�_�  F  I          G   �        ����                                                                                                                                                                                                                                                                                                                            �           �   >          >    Z �     �   �   �   �      //�   �   �   �    5�_�  G  J  H      I   �        ����                                                                                                                                                                                                                                                                                                                            �           �   >          >    Z �     �   �   �   �       �   �   �   �    5�_�  I  K          J   �        ����                                                                                                                                                                                                                                                                                                                            �           �   >          >    Z �     �   �   �   �                       �   �   �   �    5�_�  J  L          K   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �      milk_remain     > milk_req        chocolate_remain> chocolate_req   froth_remain    > froth_req    �   �   �   �      espresso_remain > espresso_req 5�_�  K  M          L   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �      != milk_remain     > milk_req        != chocolate_remain> chocolate_req   != froth_remain    > froth_req    �   �   �   �      != espresso_remain > espresso_req 5�_�  L  N          M   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �              �   �   �   �    5�_�  M  O          N   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �      logic 5�_�  N  P          O   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �      logic []5�_�  O  Q          P   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �      logic []5�_�  P  R          Q   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z ��     �   �   �   �      7logic espresso_led, milk_led, chocolate_led, froth_led;5�_�  Q  S          R   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z ��     �   �   �   �      )      milk_led, chocolate_led, froth_led;�   �   �   �      7logic espresso_led, milk_led, chocolate_led, froth_led;5�_�  R  T          S   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z ��     �   �   �   �      )      milk_led, chocolate_led, froth_led;5�_�  S  U          T   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z ��     �   �   �   �      )      milk_led, chocolate_led, froth_led;5�_�  T  V          U   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z ��     �   �   �   �            chocolate_led, froth_led;�   �   �   �      -      milk_led    , chocolate_led, froth_led;5�_�  U  W          V   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z ��     �   �   �   �            froth_led;�   �   �   �            chocolate_led, froth_led;5�_�  V  X          W   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z ��     �   �   �   �            chocolate_led, �   �   �   �            froth_led;5�_�  W  Y          X   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �      �   �   �   �            milk_led    , 5�_�  X  Z          Y   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z �     �   �   �   �      logic espresso_led, 5�_�  Y  [          Z   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �
     �   �   �   �      (assign = espresso_remain > espresso_req    (assign = milk_remain     > milk_req        (assign = chocolate_remain> chocolate_req   (assign = froth_remain    > froth_req        �   �   �   �    5�_�  Z  \          [   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      5assign espresso_led = espresso_remain > espresso_req 5�_�  [  ]          \   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      5assign milk_led     = milk_remain     > milk_req     5�_�  \  ^          ]   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      5assign chocolate_led= chocolate_remain> chocolate_req5�_�  ]  _          ^   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �     �   �   �   �      5assign froth_led    = froth_remain    > froth_req    5�_�  ^  `          _   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z �&    �   �   �   �      W            espresso_remain <= ( )? espresso_remain - espresso_req  : espresso_remain ;   W            milk_remain     <= ( )? milk_remain     - milk_req      : milk_remain     ;   W            chocolate_remain<= ( )? chocolate_remain- chocolate_req : chocolate_remain;   W            froth_remain    <= ( )? froth_remain    - froth_req     : froth_remain    ;       end�   �   �   �    5�_�  _  a          `           ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �         �       �         �    5�_�  `  b          a          ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �         �      typedef struct 5�_�  a  c          b          ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �         �      typedef struct {}5�_�  b  d          c          ����                                                                                                                                                                                                                                                                                                                                                             Z ��     �         �      typedef struct {}5�_�  c  e          d          ����                                                                                                                                                                                                                                                                                                                                                             Z �(     �         �      typedef struct {} FSM_state;5�_�  d  f          e          ����                                                                                                                                                                                                                                                                                                                                                             Z �+     �         �      typedef enum {} FSM_state;5�_�  e  g          f          ����                                                                                                                                                                                                                                                                                                                                                             Z �+     �         �      typedef enum []{} FSM_state;5�_�  f  h          g          ����                                                                                                                                                                                                                                                                                                                                                             Z �,     �         �      typedef enum []{} FSM_state;5�_�  g  i          h          ����                                                                                                                                                                                                                                                                                                                                                             Z �/     �         �      typedef enum [2:0]{} FSM_state;5�_�  h  j          i          ����                                                                                                                                                                                                                                                                                                                                                             Z �1     �         �      typedef enum [2:0]{} FSM_state;5�_�  i  k          j          ����                                                                                                                                                                                                                                                                                                                                                             Z �5     �         �      $typedef enum logic[2:0]{} FSM_state;5�_�  j  l          k          ����                                                                                                                                                                                                                                                                                                                                                             Z �c     �         �      Btypedef enum logic[2:0]{S_INPUT,S_MILK,S_CHOCO,S_FROTH} FSM_state;5�_�  k  m          l      &    ����                                                                                                                                                                                                                                                                                                                                                             Z �s     �         �      Itypedef enum logic[2:0]{S_IDLE,S_INPUT,S_MILK,S_CHOCO,S_FROTH} FSM_state;5�_�  l  n          m      ,    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �         �       �         �    5�_�  m  o          n          ����                                                                                                                                                                                                                                                                                                                                                             Z �     �         �    5�_�  n  q          o      D    ����                                                                                                                                                                                                                                                                                                                                                             Z �     �         �      Ptypedef enum logic[2:0]{S_IDLE,S_INPUT,S_ESPR,S_MILK,S_CHOCO,S_FROTH} FSM_state;5�_�  o  r  p      q          ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �+    �         �      ttypedef enum logic[2:0]{S_IDLE,S_INPUT,S_ESPR,S_MILK,S_CHOCO,S_FROTH,S_CUSTO_BASE,S_COMP_UPDATE,S_OUTPUT} FSM_state;5�_�  q  s          r   �        ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �7     �   �   �   �       �   �   �   �    5�_�  r  t          s   �   
    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �D     �   �   �   �      
always_ff@5�_�  s  u          t   �   +    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �K     �   �   �   �      ,always_ff@(posedge clk or negedge inf.rst_n)5�_�  t  v          u   �   ,    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �K     �   �   �   �      ,always_ff@(posedge clk or negedge inf.rst_n)5�_�  u  w          v   �   0    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �L     �   �   �   �          �   �   �   �    5�_�  v  x          w   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �M     �   �   �   �          �   �   �   �    5�_�  w  y          x   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �O     �   �   �   �          if5�_�  x  z          y   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �R     �   �   �   �          if(inf.rst_n)5�_�  y  {          z   �   
    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �S     �   �   �   �          if(inf.rst_n)5�_�  z  |          {   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �S     �   �   �   �          if(inf.rst_n)5�_�  {  }          |   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �T     �   �   �   �          if(inf.rst_n)5�_�  |  ~          }   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �W     �   �   �   �          if(!inf.rst_n)5�_�  }            ~   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �X     �   �   �   �              �   �   �   �    5�_�  ~  �             �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �Y     �   �   �   �    5�_�    �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �Z     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �\     �   �   �   �              �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �\     �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �^     �   �   �   �       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �n     �   �   �   �              �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �w     �   �   �           5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �x     �   �   �   �       �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �      always_comb@5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �      always_comb@()5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �      always_comb@()5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �          �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �          case5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �          case(c_state)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �              �   �   �   �    5�_�  �  �          �   �   
    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �   �   �   �              �   �   �   �    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �      !   �       �          �    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �      !   �      logic invalid = 5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �      !   �      logic invalid = ()5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �      !   �      logic invalid = ()5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z ��     �      !   �      logic invalid = (inf.)5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z ��     �      !   �      (logic invalid = (inf.select_i || supply)5�_�  �  �          �       *    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z ��     �      !   �      *logic fill_flag = (inf.select_i || supply)5�_�  �  �          �       -    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z ��     �      !   �      -logic fill_flag = (inf.select_i || supply)? 15�_�  �  �          �       7    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z ��     �       "   �       �       "   �    5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �       "   �      logic customize = 5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �       "   �      logic customize = ()5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �       "   �      logic customize = ()5�_�  �  �          �   !   1    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �.     �       "   �      1logic customize = (inf.flavor_btn == user_define)5�_�  �  �          �   !   5    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �/     �       "   �      5logic customize = (inf.flavor_btn == user_define) ? 15�_�  �  �          �   !   ?    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �K     �   !   #   �       �   !   #   �    5�_�  �  �          �   "        ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �z    �   !   "          logic in_valid  =5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z ��    �      !   �       �      !   �    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �[     �         �      ttypedef enum logic[3:0]{S_IDLE,S_INPUT,S_ESPR,S_MILK,S_CHOCO,S_FROTH,S_CUSTO_BASE,S_COMP_UPDATE,S_OUTPUT} FSM_state;5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                            !          #          V       Z �h     �       !          %// ------------ flag ----------------   8logic fill_flag = (inf.select_i || supply)? 1'b1 : 1'b0;   @logic customize = (inf.flavor_btn == user_define) ? 1'b1 : 1'b0;5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �l     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �v     �   �   �   �              S_IDLE:5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �      +        S_IDLE:(fill_flag || customize || )5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �      +        S_IDLE:(fill_flag || customize || )5�_�  �  �          �   �   8    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �      8        S_IDLE:(fill_flag || customize || required_size)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �                  �   �   �   �    5�_�  �  �          �   �   
    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �                  �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �                  if5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �                  if(customize)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �                  if(customize)5�_�  �  �          �   �   $    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �                  �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �   �   �   �                  else if5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �                  else if()5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �                  else if()5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �      @logic customize = (inf.flavor_btn == user_define) ? 1'b1 : 1'b0;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �                  if(customize)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �                  else if(fill_flag)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �                  else if(fill_flag)b5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �   �   �                      �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �%     �   �   �   �                  �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �)     �   �   �   �                  else if5�_�  �  �          �   �   !    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �0     �   �   �   �      "            else if(required_size)5�_�  �  �          �   �   "    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �2     �   �   �   �      "            else if(required_size)5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �C     �   �   �   �                  �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �F     �   �   �   �                      �   �   �   �    5�_�  �  �          �   �   
    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �L     �   �   �                 �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �e     �   �   �      5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �h     �   �   �                    �   �   �      5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �o     �   �                           �   �         5�_�  �  �          �   �   %    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �w     �   �                      �   �        5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �                      S_CHOCOLATE:5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �   �                  S_CHOCOLATE:5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �                        �           5�_�  �  �          �     !    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �                        �          5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �                            �          5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �      	                  �          5�_�  �  �          �     
    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �      	                  S_FROTH:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �      
                    �      	    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �                            �      
    5�_�  �  �          �     '    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �          5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �                        S_CUSTO_BASE:5�_�  �  �          �     
    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �                      S_FROTH:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �                    S_CUSTO_BASE:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �                 S_CUSTO_BASE:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �                 S_CUSTO_BASE:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z ��     �                        �          5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �                        S_COMP_UPDATE:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �                    S_COMP_UPDATE:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �     �            	         �          5�_�  �  �          �  	       ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �!     �    	                          5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �"     �               5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �#     �               5�_�  �  �          �      S    ����                                                                                                                                                                                                                                                                                                                            !          !          V       Z �F    �              e        {S_IDLE,S_INPUT,S_ESPR,S_MILK,S_CHOCO,S_FROTH,S_CUSTO_BASE,S_COMP_UPDATE,S_OUTPUT} FSM_state;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-I     �            5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-K    �                 5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-Q     �            5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-S    �                 5�_�  �  �  �      �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �            5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�    �                 5�_�  �  �          �            ����                                                                                                                                                                                                                                                                                                                                                             Z!-�    �                  5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �   �   �  
    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z!-�    �   �   �           5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �                 5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �        	    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�    �                 5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �        	    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �                 5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �        	    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�   " �                 5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                                                             Z!-�   $ �        	    5�_�  �  �          �   <        ����                                                                                                                                                                                                                                                                                                                                                             Z!.   % �   ;   <           5�_�  �  �          �   I        ����                                                                                                                                                                                                                                                                                                                                                             Z!.   & �   H   I           5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                             Z!.     �              logic [3:0] base;   logic [5:0] weight_size;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             Z!.     �              *logic [3:0] base; logic [5:0] weight_size;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             Z!.   ' �              )logic [3:0] base;logic [5:0] weight_size;5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                                                             Z!.+     �       "        always_comb   begin: base_selector5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                                                             Z!.,   ( �       #         always_comb begin: base_selector5�_�  �  �          �   =        ����                                                                                                                                                                                                                                                                                                                                                             Z!.7   ) �   =   ?  	      // �   =   ?      5�_�  �  �          �   9        ����                                                                                                                                                                                                                                                                                                                                                             Z!.J     �   9   ;  	    5�_�  �  �          �   :        ����                                                                                                                                                                                                                                                                                                                                                             Z!.K   * �   9   :           5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             Z!9     �        	      b        {S_IDLE,S_INPUT,S_ESPR,S_MILK,S_CHOCO,S_FROTH,S_CUSTO_BASE,S_COMP_UPDAT_OUTPUT} FSM_state;5�_�  �  �          �   C       ����                                                                                                                                                                                                                                                                                                                                                             Z!9     �   B   D  	      %    else if(n_state == S_INPUT)begin 5�_�  �  �          �   O       ����                                                                                                                                                                                                                                                                                                                                                             Z!9J     �   N   P  	      &    else if(n_state == S_INPUT) begin 5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                                                             Z!9z   + �   <   >  	      :// -------------------  S_INPUT --------------------------5�_�  �  �          �   C   $    ����                                                                                                                                                                                                                                                                                                                                                             Z!=      �   B   D  	      +    else if(n_state == S_GENERAL_REQ)begin 5�_�  �  �          �   O   $    ����                                                                                                                                                                                                                                                                                                                                                             Z!=M     �   N   P  	      ,    else if(n_state == S_GENERAL_REQ) begin 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!=�     �   �   �  	                  S_ESPRESSO:begin5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!=�     �   �   �  	                  S_ESPR:begin5�_�  �  �          �   O   9    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!=�     �   N   P  	      A    else if(n_state == S_GENERAL_REQ || n_state == S_ESPR) begin 5�_�  �  �          �   C   9    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!=�     �   B   D  	      @    else if(n_state == S_GENERAL_REQ || n_state == S_ESPR)begin 5�_�  �             �      $    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!=�     �        	      h        {S_IDLE,S_GENERAL_REQ,S_ESPR,S_MILK,S_CHOCO,S_FROTH,S_CUSTO_BASE,S_COMP_UPDAT_OUTPUT} FSM_state;5�_�  �                �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>!     �   �   �  	    5�_�                  �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>0     �   �   �  
       5�_�                 �   
    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>4     �   �   �  
      
always_ff@5�_�                 �   !    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>B     �   �   �  
      "always_ff@(posedge clk or negedge)5�_�                 �   !    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>F     �   �   �  
      "always_ff@(posedge clk or negedge)5�_�                 �   ,    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>K     �   �   �  
      ,always_ff@(posedge clk or negedge inf.rst_n)5�_�                 �   0    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>L     �   �   �            �   �   �  
    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>M     �   �   �            �   �   �      5�_�    	             �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>O     �   �   �            if5�_�    
          	   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>U     �   �   �            if(! inf.rst_n)5�_�  	            
   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>U     �   �   �            if(! inf.rst_n)5�_�  
               �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>W     �   �   �                �   �   �      5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>X     �   �   �                �   �   �      5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>a     �   �   �                sum_weight <= 5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>c     �   �   �                sum_weight <= 'b0;'5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>d     �   �   �                sum_weight <= 'b0;'5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>e     �   �   �            �   �   �      5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>g     �   �   �            else if5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>l     �   �   �            else if(S_IDLE)5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>r     �   �   �            else if(S_IDLE)5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>y     �   �   �            else if(n_state == S_IDLE)5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>{     �   �   �      5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if(n_state == S_IDLE)5�_�                 �   "    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �                �   �   �      5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �                �   �   �      5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �                sum_weight <= 5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �                sum_weight <= 'b0'5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �                sum_weight <= 'b0'5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            �   �   �      5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if5�_�                  �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            �   �   �      5�_�    !            �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if5�_�     "          !   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if5�_�  !  #          "   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if5�_�  "  $          #   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if()5�_�  #  %          $   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if()5�_�  $  &          %   �   A    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?;     �   �   �        B    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state)5�_�  %  '          &   �   B    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?H     �   �   �        U    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state || S_CHOCOLATE || )5�_�  &  (          '   �   B    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?H     �   �   �        T    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state | S_CHOCOLATE || )5�_�  '  )          (   �   B    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?J     �   �   �        S    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state  S_CHOCOLATE || )5�_�  (  *          )   �   F    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?K     �   �   �        U    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state == S_CHOCOLATE || )5�_�  )  +          *   �   T    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?N     �   �   �        U    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state == S_CHOCOLATE || )5�_�  *  ,          +   �   b    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?Y     �   �   �        c    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state == S_CHOCOLATE || n_state == S_C)5�_�  +  -          ,   �   f    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?c     �   �   �        l    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state == S_CHOCOLATE || n_state == S_CUSTO_BASE)5�_�  ,  .          -   �   :    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?k     �   �   �        m    else if(n_state == S_ESPRESSO || n_state == S_MILK || n_state == S_CHOCOLATE || n_state == S_CUSTOM_BASE)5�_�  -  /          .   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?r   , �   �   �                    �   �   �      5�_�  .  0          /   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?�     �   �   �          (    else if(flavor_btn_r == user_define)5�_�  /  1          0   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?�     �   �   �                �   �   �      5�_�  0  2          1   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?�     �   �   �                �   �   �      5�_�  1  3          2   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?�     �   �   �           5�_�  2  4          3   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?�     �   �   �      5�_�  3  5          4   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?�     �   �   �        Xassign sum_weight = (espresso_weight + milk_weight) + (chocolate_weight + froth_weight);5�_�  4  6          5   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!?�     �   �   �        Xassign sum_weight = (espresso_weight + milk_weight) + (chocolate_weight + froth_weight);5�_�  5  7          6   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A     �   �   �      5�_�  6  8          7   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A     �   �   �        7assign user_define_base = ingredient_base / sum_weight;5�_�  7  9          8   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A     �   �   �        7assign user_define_base = ingredient_base / sum_weight;5�_�  8  :          9   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A     �   �   �        //�   �   �      5�_�  9  ;          :   �   
    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A#     �   �   �        
always_ff@5�_�  :  <          ;   �   +    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A(     �   �   �        ,always_ff@(posedge clk or negedge inf.rst_n)5�_�  ;  =          <   �   ,    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A(     �   �   �        ,always_ff@(posedge clk or negedge inf.rst_n)5�_�  <  >          =   �   0    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A)     �   �   �            �   �   �      5�_�  =  ?          >   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A.     �   �   �              endk5�_�  >  @          ?   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A/     �   �   �            �   �   �      5�_�  ?  A          @   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A1     �   �   �            �   �   �      5�_�  @  B          A   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A2     �   �   �            if5�_�  A  C          B   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A5     �   �   �            if(!inf.rst_n)5�_�  B  D          C   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A5     �   �   �            if(!inf.rst_n)5�_�  C  E          D   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A6     �   �   �      �   �   �      5�_�  D  F          E   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A7     �   �   �            endk5�_�  E  G          F   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A9     �   �   �            if(!inf.rst_n)begom5�_�  F  H          G   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A:     �   �   �            if(!inf.rst_n)bego5�_�  G  I          H   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A<     �   �   �                �   �   �      5�_�  H  J          I   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AC     �   �   �            end5�_�  I  K          J   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AD     �   �   �            �   �   �      5�_�  J  L          K   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AF     �   �   �                �   �   �      5�_�  K  M          L   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AG     �   �   �      5�_�  L  N          M   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AH     �   �   �                 5�_�  M  O          N   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AR     �   �   �                 user_define_base <= 5�_�  N  P          O   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AS     �   �   �                  user_define_base <= 'b0'5�_�  O  Q          P   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!AS     �   �   �                  user_define_base <= 'b0'5�_�  P  R          Q   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A[     �   �   �  !              �   �   �       5�_�  Q  S          R   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!Ah     �   �   �  !              user_define_base <= 5�_�  R  T          S   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!Ah     �   �   �  !              user_define_base <= ()5�_�  S  V          T   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!Az     �   �   �  !              user_define_base <= ()5�_�  T  W  U      V   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A�     �   �   �  !      6        user_define_base <= (c_state == S_CUSTOM_BASE)�   �   �  !    5�_�  V  X          W   �   8    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A�     �   �   �  !      8        user_define_base <= (c_state == S_CUSTOM_BASE)//5�_�  W  Y          X   �   V    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A�     �   �   �  !      V        user_define_base <= (c_state == S_CUSTOM_BASE) ? ingredient_base/sum_weight : 5�_�  X  Z          Y   �   Z    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A�     �   �   �  !      Z        user_define_base <= (c_state == S_CUSTOM_BASE) ? ingredient_base/sum_weight : user5�_�  Y  [          Z   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A�     �   �   �           5�_�  Z  \          [   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!B*     �   �   �           5�_�  [  ]          \   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!BX     �   �   �        6assign milk_led     = milk_remain     > milk_req     ;   6assign chocolate_led= chocolate_remain> chocolate_req;   6assign froth_led    = froth_remain    > froth_req    ;�   �   �        6assign espresso_led = espresso_remain > espresso_req ;5�_�  \  ^          ]   �   6    ����                                                                                                                                                                                                                                                                                                                            �   6       �   6          6    Z!B]     �   �   �        7assign espresso_led = (espresso_remain > espresso_req ;5�_�  ]  _          ^   �   ;    ����                                                                                                                                                                                                                                                                                                                            �   6       �   6          6    Z!Ba     �   �   �        7assign milk_led     = (milk_remain     > milk_req     ;   7assign chocolate_led= (chocolate_remain> chocolate_req;   7assign froth_led    = (froth_remain    > froth_req    ;�   �   �        <assign espresso_led = (espresso_remain > espresso_req ) ? 1;5�_�  ^  `          _   �   #    ����                                                                                                                                                                                                                                                                                                                            �   6       �   6          6    Z!B|     �   �   �        8logic fill_flag = (inf.select_i || supply)? 1'b1 : 1'b0;5�_�  _  a          `   �   "    ����                                                                                                                                                                                                                                                                                                                            �   "       �   <          <    Z!B�     �   �   �        dlogic [9:0]  ingredient_basis  = (flavor_btn_r == user_define) ? user_define_base : ingredient_base;5�_�  `  b          a   �   "    ����                                                                                                                                                                                                                                                                                                                            �   "       �   <          <    Z!B�   - �   �   �        Ilogic [9:0]  ingredient_basis  = () ? user_define_base : ingredient_base;5�_�  a  c          b   �        ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�     �   �   �          %// ------------ flag ----------------   <logic fill_flag = (inf.select_i || inf.supply)? 1'b1 : 1'b0;   Elogic customize_flag = (inf.flavor_btn == user_define) ? 1'b1 : 1'b0;5�_�  b  d          c           ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�     �            �            5�_�  c  e          d           ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�   . �      !          �             5�_�  d  f          e         ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�     �                         S_FROTH:5�_�  e  g          f         ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�     �              '                n_state = S_CUSTO_BASE;5�_�  f  h          g         ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�     �            "                n_state = S_FROTH;5�_�  g  i          h         ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�     �                            n_state = S;5�_�  h  j          i         ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�     �                  S_CUSTO_BASE:5�_�  i  k          j   "   G    ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!B�   / �   !   #        l        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_FROTH,S_CUSTO_BASE,S_COMP_UPDAT_OUTPUT} FSM_state;5�_�  j  l          k   �       ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!C1     �   �   �                    S_FROTH:begin5�_�  k  m          l   q       ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!C=     �   q   s                         �   q   s      5�_�  l  n          m   r       ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!C>     �   q   s                         if5�_�  m  o          n   r   !    ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!CB     �   q   s         "                if(customize_flag)5�_�  n  p          o   r   "    ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!CD     �   q   s         "                if(customize_flag)5�_�  o  q          p   r   &    ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!CF     �   r   t  !                          �   r   t       5�_�  p  r          q   r       ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!CH     �   r   t  !    5�_�  q  s          r   t       ����                                                                                                                                                                                                                                                                                                                            �   $       �   /       V   /    Z!CI     �   t   v  #                      �   t   v  "    5�_�  r  t          s   �       ����                                                                                                                                                                                                                                                                                                                               $          /       V   /    Z!CM     �   �   �  $                      �   �   �  #    5�_�  s  u          t   v       ����                                                                                                                                                                                                                                                                                                                            v          �                 Z!CR     �   v   �  $                           latte: begin   0                        espresso_weight <= 3'd2;   0                        milk_weight      <=3'd1;   0                        chocolate_weight <=3'd0;   0                        froth_weight     <=3'd2;                       end   $                    cappuccino:begin   0                        espresso_weight <= 3'd2;   0                        milk_weight      <=3'd1;   0                        chocolate_weight <=3'd0;   0                        froth_weight     <=3'd1;                       end                        mocha: begin   0                        espresso_weight <= 3'd1;   0                        milk_weight      <=3'd1;   0                        chocolate_weight <=3'd1;   0                        froth_weight     <=3'd0;                       end                       default:   0                        espresso_weight <= 3'd0;   0                        milk_weight      <=3'd0;   0                        chocolate_weight <=3'd0;   0                        froth_weight     <=3'd0;                   endcase�   u   w  $                       case(flavor_btn)5�_�  t  w          u   �       ����                                                                                                                                                                                                                                                                                                                            v          �                 Z!CV     �   �   �  $                  end5�_�  u  y  v      w   r       ����                                                                                                                                                                                                                                                                                                                            x          {   +          +    Z!Ch     �   r   v  %                          �   r   t  $    5�_�  w  z  x      y   s        ����                                                                                                                                                                                                                                                                                                                            {          ~   +          +    Z!Ck     �   r   x  '                                      end�   s   t  '    5�_�  y  {          z   s        ����                                                                                                                                                                                                                                                                                                                            s           v                   Z!Cn     �   s   w  '      milk_weight        chocolate_weight   froth_weight    �   r   t  '      espresso_weight 5�_�  z  |          {   s   ,    ����                                                                                                                                                                                                                                                                                                                            s           v                   Z!Cr     �   r   t  '      ,                            espresso_weight 5�_�  {  }          |   s   ,    ����                                                                                                                                                                                                                                                                                                                            s   ,       v   ,          ,    Z!Cv     �   s   w  '      ,                            milk_weight        ,                            chocolate_weight   ,                            froth_weight    �   r   t  '      -                            espresso_weight  5�_�  |  ~          }   s   -    ����                                                                                                                                                                                                                                                                                                                            s   -       v   -          -    Z!Cy     �   r   w  '      0                            espresso_weight < =    /                            milk_weight     < =   /                            chocolate_weight< =   /                            froth_weight    < =5�_�  }            ~   s   .    ����                                                                                                                                                                                                                                                                                                                            s          v   +          +    Z!C     �   r   x  '      /                            espresso_weight <=    .                            milk_weight     <=   .                            chocolate_weight<=   .                            froth_weight    <=                   end�   s   t  '    5�_�  ~  �             s   ?    ����                                                                                                                                                                                                                                                                                                                            s   >       v   >          >    Z!C�   0 �   s   w  '      ?                            milk_weight     <= milk_weight        ?                            chocolate_weight<= chocolate_weight   ?                            froth_weight    <= froth_weight    �   r   t  '      ?                            espresso_weight <= espresso_weight 5�_�    �          �   y   #    ����                                                                                                                                                                                                                                                                                                                            s   >       v   >          >    Z!C�     �   x   z  '      $                    case(flavor_btn)5�_�  �  �          �   r       ����                                                                                                                                                                                                                                                                                                                            s   >       v   >          >    Z!C�     �   q   r          '                if(customize_flag)begin5�_�  �  �          �   r        ����                                                                                                                                                                                                                                                                                                                            r          u          V       Z!C�     �   q   r          @                            espresso_weight <= espresso_weight ;   @                            milk_weight     <= milk_weight     ;   @                            chocolate_weight<= chocolate_weight;   @                            froth_weight    <= froth_weight    ;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            r          r          V       Z!C�     �   �   �  "    �   �   �  "    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            r          r          V       Z!C�     �   �   �  '                              �   �   �  &    5�_�  �  �          �   �   (    ����                                                                                                                                                                                                                                                                                                                            r          r          V       Z!C�     �   �   �  (                                  �   �   �  '    5�_�  �  �          �   r       ����                                                                                                                                                                                                                                                                                                                            r          r          V       Z!C�     �   q   r                          end5�_�  �  �          �   r       ����                                                                                                                                                                                                                                                                                                                            r          r          V       Z!C�     �   q   r                          else begin5�_�  �  �          �   �   ,    ����                                                                                                                                                                                                                                                                                                                            r          r          V       Z!C�   1 �      �  &      4                            espresso_weight <= 3'd1;5�_�  �  �  �      �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z!DG     �   �   �  &          else begin5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z!DI     �   �   �  &          else if begin5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                            �           �                   Z!DP     �   �   �  &      1    else if(c_state == S_COMP_UPDAT_OUTPUT) begin5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �           �                   Z!DR     �       '          �       &    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �           �                   Z!DT     �      (              �      '    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �           �                   Z!DU     �      (    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!D^     �      *              �      )    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!D`     �      ,       5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!Da     �      ,                                     end�      ,    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                                     Z!Dg     �      ,                  milk_remain                    chocolate_remain               froth_remain    �      ,                  espresso_remain 5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                                     Z!Dj     �      ,                   espresso_remain  <=                 milk_remain      <=                 chocolate_remain <=                 froth_remain     <=        end�      ,    5�_�  �  �          �     /    ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!Dm     �      ,      0            milk_remain      <=milk_remain         0            chocolate_remain <=chocolate_remain    0            froth_remain     <=froth_remain     �      ,      0            espresso_remain  <=espresso_remain  5�_�  �  �          �     /    ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!Dq   4 �      ,      1            espresso_remain  <=espresso_remain l    1            milk_remain      <=milk_remain     l    1            chocolate_remain <=chocolate_remainl    1            froth_remain     <=froth_remain    l 5�_�  �  �          �   "   8    ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!H�     �   !   #  ,      m        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_FROTH,S_CUSTOM_BASE,S_COMP_UPDAT_OUTPUT} FSM_state;5�_�  �  �          �   "   8    ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!H�   5 �   !   #  ,      f        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,,S_CUSTOM_BASE,S_COMP_UPDAT_OUTPUT} FSM_state;5�_�  �  �          �            ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!H�   6 �                  5�_�  �  �          �   !   Y    ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!I   7 �       "  +      e        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_CUSTOM_BASE,S_COMP_UPDAT_OUTPUT} FSM_state;5�_�  �  �  �      �   �   #    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�     �   �   �  +      1    else if(c_state == S_COMP_UPDAT_OUTPUT) begin5�_�  �  �          �   �   #    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�     �   �   �  +      )    else if(c_state == S_COMP_UPDAT begin5�_�  �  �          �   !   R    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�     �       "  +      l        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_CUSTOM_BASE,S_COMP_UPDAT_OUTPUT,S_FILL} FSM_state;5�_�  �  �          �   !   S    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�     �       "  +      l        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_CUSTOM_BASE,S_COMP_UPDATeOUTPUT,S_FILL} FSM_state;5�_�  �  �          �   !   R    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�     �       "  +      f        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_CUSTOM_BASE,S_COMP_UPDATe,S_FILL} FSM_state;5�_�  �  �          �   !   R    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�   8 �       "  +      e        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_CUSTOM_BASE,S_COMP_UPDAT,S_FILL} FSM_state;5�_�  �  �          �  %       ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�     �  $  &  +      (                n_state = S_COMP_UPDATE;5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!I�     �  %  '  +           S_COMP_UPDATE:5�_�  �  �          �  %       ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J     �  %  '  ,                  �  %  '  +    5�_�  �  �          �  &       ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J   9 �  &  (  -      
          �  &  (  ,    5�_�  �  �          �  )        ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �  )  +  .                  �  )  +  -    5�_�  �  �          �  *       ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�   : �  *  ,  /                      �  *  ,  .    5�_�  �  �          �      	    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �   �    /          else begin5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �   �    /          else ifbegin5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �       0              �       /    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �       0    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �      2          �      1    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �      2    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �       4              �       3    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �       4                  case5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!J�     �       4                  case()5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K      �   �    4      #    else if(c_state == S_FILL)begin5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K     �   �   �  4      +    else if(c_state == S_COMP_UPDATE) begin5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!Kp     �       4                  case()5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!Ku     �      5                      �      4    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!Kw     �      6                      �      5    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K     �      7                      �      6    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      7                      latte5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      7                      cappuccino5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      8                      �      7    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      8    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �                              latte:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �                              cappuccino:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �                              mocha:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �       6                  case(supply)5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      7                      �      6    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      8                          �      7    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      9                      �      8    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :                      �      9    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :                      espresso:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :                      milk:5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :                      chocolate:5�_�  �  �          �     )    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :      *                chocolate:chocolate      <5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :      +                chocolate:chocolate       <5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :                      froth:5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!K�     �      :       5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L     �      :      F                espresso: espresso_remain <= espresso_remain + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L     �      :      K                espresso:begin espresso_remain <= espresso_remain + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L     �      <                          �      ;    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L     �      =                          �      <    5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L     �      >                          �      =    5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L     �      >      ,                    milk            <= milk;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L     �      >      3                    milk            <= milk_remain;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L      �      >      ;                    milk_remaink            <= milk_remain;5�_�  �  �          �     $    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L#     �      >      :                    milk_remain            <= milk_remain;5�_�  �  �          �     #    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L&     �      >      7                    chocolate       M= chocolate_remain5�_�  �  �          �     #    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L'     �      >      6                    chocolate      M= chocolate_remain5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L)     �      >      5                    chocolate      = chocolate_remain5�_�  �  �          �     %    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L,     �      >      =                    chocolate_remaine      = chocolate_remain5�_�  �  �          �     %    ����                                                                                                                                                                                                                                                                                                                            �   #       �   *          *    Z!L-     �      >      7                    chocolate_remaine= chocolate_remain5�_�  �  �          �     $    ����                                                                                                                                                                                                                                                                                                                              $         $          $    Z!L1     �      >      3                    milk_remain     <= milk_remain;�      >      @                    espresso_remain <= espresso_remain + supply;5�_�  �  �          �     $    ����                                                                                                                                                                                                                                                                                                                              $         $          $    Z!L3     �      ?                          �      >    5�_�  �  �          �     &    ����                                                                                                                                                                                                                                                                                                                              $         $          $    Z!L:     �      ?      (                    froth_remain        5�_�  �  �          �     9    ����                                                                                                                                                                                                                                                                                                                              $         $          $    Z!LB     �      ?      9                    chocolate_remaine <= chocolate_remain5�_�  �  �          �     $    ����                                                                                                                                                                                                                                                                                                                              $         $          $    Z!LE     �      ?      :                    chocolate_remaine <= chocolate_remain;5�_�  �  �          �     %    ����                                                                                                                                                                                                                                                                                                                              $         $          $    Z!LF   ; �      ?      9                    chocolate_remain <= chocolate_remain;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!LS     �    	  ?      F                milk:     milk            <= milk            + supply;5�_�  �  �          �     &    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!LU     �    	  ?      M                milk:     milk_remain            <= milk            + supply;5�_�  �  �          �     .    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!LX     �    	  ?      B                milk:     milk_remain <= milk            + supply;5�_�  �  �          �     8    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L\     �    	  ?      H                milk:     milk_remain <= milk_remain           + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!Lc     �    	  ?      A                milk:     milk_remain <= milk_remain    + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!Ld     �    
  ?    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!Lg     �    
  @      F                milk:begin     milk_remain <= milk_remain    + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!Li     �    
  B                      �    
  A    5�_�  �  �          �  
        ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!Lu     �  	    B      ;                    milk_remain <= milk_remain    + supply;5�_�  �  �          �  
        ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!Lz     �  
    B    �  
    B    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L|     �      E                          �      D    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �               5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      D      F                chocolate:chocolate       <= chocolate       + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      D      K                chocolate:beginchocolate       <= chocolate       + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      E    �      E    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      F    �      F    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      G      @                    chocolate       <= chocolate       + supply;5�_�  �  �          �     &    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      G      G                    chocolate_remain       <= chocolate       + supply;5�_�  �  �          �     2    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      G      B                    chocolate_remain  <= chocolate       + supply;5�_�  �  �          �     <    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      G      I                    chocolate_remain  <= chocolate_remain       + supply;5�_�  �  �          �     :    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      G      E                    chocolate_remain  <= chocolate_remain   + supply;5�_�  �  �          �     B    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      G    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      H    �      H    5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      J                          �      I    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �               5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      I      F                froth:    froth           <= froth           + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      I      K                froth:begin    froth           <= froth           + supply;5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      J      A                     froth           <= froth           + supply;5�_�  �  �          �     &    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      J      D                     froth_remain       <= froth           + supply;5�_�  �  �          �     .    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      J      B                     froth_remain     <= froth           + supply;5�_�  �  �          �     9    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      J      I                     froth_remain     <= froth_remain           + supply;5�_�  �            �     9    ����                                                                                                                                                                                                                                                                                                                              %         %       V   %    Z!L�     �      J      B                     froth_remain     <= froth_remain    + supply;5�_�  �                     ����                                                                                                                                                                                                                                                                                                                              8         5       V   9    Z!L�     �      J    �      J    5�_�                       ����                                                                                                                                                                                                                                                                                                                              8         5       V   9    Z!L�     �      L      C                     froth_remain     <= froth_remain     + supply;5�_�                       ����                                                                                                                                                                                                                                                                                                                              8         5       V   9    Z!L�     �      L    �      L    5�_�                        ����                                                                                                                                                                                                                                                                                                                                              V       Z!L�     �      M    �      M    5�_�                       ����                                                                                                                                                                                                                                                                                                                                              V       Z!L�     �      P                      default:5�_�                       ����                                                                                                                                                                                                                                                                                                                                              V       Z!L�     �      P      !                    default:begin5�_�                       ����                                                                                                                                                                                                                                                                                                                                              V       Z!L�     �      Q                          �      P    5�_�    	                   ����                                                                                                                                                                                                                                                                                                                                              V       Z!L�     �      Q    �      Q    5�_�    
          	           ����                                                                                                                                                                                                                                                                                                                                              V       Z!L�     �                5�_�  	            
           ����                                                                                                                                                                                                                                                                                                                                              V       Z!L�     �                5�_�  
              J       ����                                                                                                                                                                                                                                                                                                                                              V       Z!M     �  J  L  Q                  �  J  L  P    5�_�                K       ����                                                                                                                                                                                                                                                                                                                                              V       Z!M   = �  K  M  R                      �  K  M  Q    5�_�                P        ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  P  S  S       �  P  R  R    5�_�                R   
    ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  Q  S  T      
always_ff@5�_�                R   +    ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  Q  S  T      ,always_ff@(posedge clk or negedge inf.rst_n)5�_�                R   ,    ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  Q  S  T      ,always_ff@(posedge clk or negedge inf.rst_n)5�_�                R   0    ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  R  T  U          �  R  T  T    5�_�                R       ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  R  T  V          �  R  T  U    5�_�                S       ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  R  T  V          if5�_�                S       ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  R  T  V          if(!inf.rst_n)5�_�                S       ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  R  T  V          if(!inf.rst_n)5�_�                S       ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  S  U  W              �  S  U  V    5�_�                S       ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  S  U  W    5�_�                U       ����                                                                                                                                                                                                                                                                                                                                              V       Z!O�     �  U  W  Y          �  U  W  X    5�_�                V       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P      �  V  X  Z              �  V  X  Y    5�_�                W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  V  X  Z              endk5�_�                V   
    ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  V  X  [              �  V  X  Z    5�_�                X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  W  Y  [              end5�_�                V       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  V  X  \              �  V  X  [    5�_�                W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  V  X  \              case5�_�                 W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  V  X  \              case(n_state)5�_�    !             W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  W  Y  ]                  �  W  Y  \    5�_�     "          !  W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  W  Y  ]    5�_�  !  #          "  Z       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P     �  Y  Z                  5�_�  "  $          #  P       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P`     �  P  T  ]    �  P  Q  ]    5�_�  #  %          $  P       ����                                                                                                                                                                                                                                                                                                                                              V       Z!Pb     �  P  R  a       �  P  R  `    5�_�  $  &          %  Q       ����                                                                                                                                                                                                                                                                                                                                              V       Z!Pf     �  P  R  a      /*           output  out_valid,5�_�  %  '          &  R       ����                                                                                                                                                                                                                                                                                                                                              V       Z!Pg     �  Q  S  `              output	window,5�_�  &  (          '  S       ����                                                                                                                                                                                                                                                                                                                                              V       Z!Ph     �  R  T  `              output	flavor_out5�_�  '  )          (  S       ����                                                                                                                                                                                                                                                                                                                                              V       Z!Pj     �  R  T  `         output	flavor_out5�_�  (  *          )  V       ����                                                                                                                                                                                                                                                                                                                                              V       Z!Pw     �  V  X  a              �  V  X  `    5�_�  )  +          *  W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!Pz     �  V  X  a              out_valid <= 15�_�  *  ,          +  W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P|     �  W  Y  b              �  W  Y  a    5�_�  +  -          ,  W       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  V  X  b              out_valid <= 1'b0;5�_�  ,  .          -  X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  W  Y  b              window5�_�  -  /          .  X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  W  Y  b              inf.window5�_�  .  0          /  X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  X  Z  c              �  X  Z  b    5�_�  /  1          0  X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  W  Y  c              inf.window 5�_�  0  2          1  X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  W  Y  c              inf.window    <=5�_�  1  3          2  X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  W  Y  c              inf.window    <= 5�_�  2  4          3  X       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  X  Z  c    �  X  Y  c    5�_�  3  5          4  Y       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  Y  [  d    �  Y  Z  d    5�_�  4  6          5  Z       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  Z  \  e    �  Z  [  e    5�_�  5  7          6  Y       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  X  Z  f      "        inf.window.espresso    <= 5�_�  6  8          7  Z       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�     �  Y  [  f      "        inf.window.espresso    <= 5�_�  7  ;          8  [       ����                                                                                                                                                                                                                                                                                                                                              V       Z!P�   ? �  Z  \  f      "        inf.window.espresso    <= 5�_�  8  <  9      ;   �        ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �   �   �          #            espresso_remain <= 'b0;5�_�  ;  =          <   �        ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �   �   �          d            espresso_remain <= (espresso_led  )? espresso_remain - espresso_req  : espresso_remain ;5�_�  <  >          =          ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �              B                    espresso_remain   <= espresso_remain + supply;5�_�  =  ?          >  	        ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �    
          9                    espresso_remain   <= espresso_remain;5�_�  >  @          ?          ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �              9                    espresso_remain   <= espresso_remain;5�_�  ?  A          @          ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �              9                    espresso_remain   <= espresso_remain;5�_�  @  B          A          ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �              9                    espresso_remain   <= espresso_remain;5�_�  A  C          B  "        ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!R�     �  !  #          1            espresso_remain  <=espresso_remain ; 5�_�  B  D          C   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!R�     �   �   �          logic [9:0] espresso_remain,               milk_remain,                   chocolate_remain,               froth_remain;    5�_�  C  E          D   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!R�     �   �   �  b      Fassign espresso_led = (espresso_remain > espresso_req ) ? 1'b1 : 1'b0;5�_�  D  F          E   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �   �   �          Fassign milk_led     = (milk_remain     > milk_req     ) ? 1'b1 : 1'b0;5�_�  E  G          F   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �   �   �          #            milk_remain     <= 'b0;5�_�  F  H          G   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �   �   �          d            milk_remain     <= (milk_led      )? milk_remain     - milk_req      : milk_remain     ;5�_�  G  I          H           ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �   �            5                    milk_remain       <= milk_remain;5�_�  H  J          I          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �              A                    milk_remain       <= milk_remain    + supply;5�_�  I  K          J          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �              5                    milk_remain       <= milk_remain;5�_�  J  L          K          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �              5                    milk_remain       <= milk_remain;5�_�  K  M          L          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �              5                    milk_remain       <= milk_remain;5�_�  L  N          M          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S     �               1            milk_remain      <=milk_remain     ; 5�_�  M  O          N   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S=     �   �   �          Fassign chocolate_led= (chocolate_remain> chocolate_req) ? 1'b1 : 1'b0;5�_�  N  P          O   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S?     �   �   �          #            chocolate_remain<= 'b0;5�_�  O  Q          P   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S@     �   �   �          d            chocolate_remain<= (chocolate_led )? chocolate_remain- chocolate_req : chocolate_remain;5�_�  P  R          Q          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SA     �               :                    chocolate_remain  <= chocolate_remain;5�_�  Q  S          R          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SB     �              :                    chocolate_remain  <= chocolate_remain;5�_�  R  T          S          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SC     �              C                    chocolate_remain  <= chocolate_remain + supply;5�_�  S  U          T          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SD     �              :                    chocolate_remain  <= chocolate_remain;5�_�  T  V          U          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SE     �              :                    chocolate_remain  <= chocolate_remain;5�_�  U  W          V           ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SF     �    !          1            chocolate_remain <=chocolate_remain; 5�_�  V  X          W   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SU     �   �   �          Fassign froth_led    = (froth_remain    > froth_req    ) ? 1'b1 : 1'b0;5�_�  W  Y          X   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SU     �   �   �          #            froth_remain    <= 'b0;5�_�  X  Z          Y   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SV     �   �   �          d            froth_remain    <= (froth_led     )? froth_remain    - froth_req     : froth_remain    ;5�_�  Y  [          Z          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SW     �              8                    froth_remain      <= froth_remain;  5�_�  Z  \          [          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SX     �    	          8                    froth_remain      <= froth_remain;  5�_�  [  ]          \          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SY     �              8                    froth_remain      <= froth_remain;  5�_�  \  ^          ]          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!SZ     �              B                    froth_remain     <= froth_remain     + supply;5�_�  ]  _          ^          ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S[     �              8                    froth_remain      <= froth_remain;  5�_�  ^  `          _  !        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!S\     �     "          1            froth_remain     <=froth_remain    ; 5�_�  _  a          `   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U     �   �   �                froth_led    ;5�_�  `  b          a   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U     �   �   �          Rassign froth_led    = (inf.window.froth.monitor    > froth_req    ) ? 1'b1 : 1'b0;5�_�  a  c          b   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U     �   �   �          �            inf.window.froth.monitor    <= (froth_led     )? inf.window.froth.monitor    - froth_req     : inf.window.froth.monitor    ;5�_�  b  d          c   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U     �   �   �                chocolate_led, 5�_�  c  e          d   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U     �   �   �          Rassign chocolate_led= (inf.window.chocolate.monitor> chocolate_req) ? 1'b1 : 1'b0;5�_�  d  f          e   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U     �   �   �          �            inf.window.chocolate.monitor<= (chocolate_led )? inf.window.chocolate.monitor- chocolate_req : inf.window.chocolate.monitor;5�_�  e  g          f   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U1     �   �   �                milk_led     , 5�_�  f  h          g   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U1     �   �   �          Rassign milk_led     = (inf.window.milk.monitor     > milk_req     ) ? 1'b1 : 1'b0;5�_�  g  i          h   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U2     �   �   �          �            inf.window.milk.monitor     <= (milk_led      )? inf.window.milk.monitor     - milk_req      : inf.window.milk.monitor     ;5�_�  h  j          i   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!U@     �   �   �          logic espresso_led , 5�_�  i  k          j   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!UC     �   �   �          Rassign espresso_led = (inf.window.espresso.monitor > espresso_req ) ? 1'b1 : 1'b0;5�_�  j  l          k   �        ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!UD     �   �   �          �            inf.window.espresso.monitor <= (espresso_led  )? inf.window.espresso.monitor - espresso_req  : inf.window.espresso.monitor ;5�_�  k  m          l   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!UJ     �   �   �           logic inf.window.espresso.led ,           inf.window.milk.led     ,           inf.window.chocolate.led,          inf.window.froth.led    ;5�_�  l  n          m   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!UK     �   �   �           5�_�  m  o          n     1    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z!U^   @ �      ]      Z                    inf.window.froth.monitor     <= inf.window.froth.monitor     + supply;5�_�  n  p          o  O        ����                                                                                                                                                                                                                                                                                                                           O   !      S          V   1    Z!Uo     �  N  O          "        inf.window.espresso    <=    "        inf.window.milk        <=    "        inf.window.chocolate   <=    "        inf.window.froth       <=            flavor_out    <= none;5�_�  o  q          p  O        ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!Uo     �  N  O           5�_�  p  r          q  Q       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!Ut     �  P  R  W              case(n_state)5�_�  q  s          r  Q   ;    ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  P  R  W      ;        case(n_state == S_COMP_UPDATE || n_state == S_FILL)5�_�  r  t          s  Q   ;    ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  P  R  W      ?        case(n_state == S_COMP_UPDATE || n_state == S_FILL)begi5�_�  s  u          t  Q       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  P  R  W      ;        case(n_state == S_COMP_UPDATE || n_state == S_FILL)5�_�  t  v          u  P   	    ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  O  Q  W          else begin5�_�  u  w          v  P   	    ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  O  Q  W      	    else 5�_�  v  x          w  P   
    ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  O  Q  W          else if   7        (n_state == S_COMP_UPDATE || n_state == S_FILL)5�_�  w  y          x  R       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  Q  R                  endcase5�_�  x  z          y  R       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  Q  R              end5�_�  y  {          z  P       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  P  R  U              �  P  R  T    5�_�  z  |          {  Q       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  P  R  U              inf.out_valid <= 15�_�  {  }          |  Q       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  Q  S  V          �  Q  S  U    5�_�  |  ~          }  R       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  R  T  W              �  R  T  V    5�_�  }            ~  S       ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  R  T  W              inf.out_valid <= 15�_�  ~  �            T        ����                                                                                                                                                                                                                                                                                                                           O   !      O          V   1    Z!U�     �  S  T           5�_�    �  �      �  H        ����                                                                                                                                                                                                                                                                                                                           H          I           V        Z!U�     �  G  H          /* output  out_valid,      output	window,5�_�  �  �          �  H       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!U�     �  G  H             output	flavor_out*/5�_�  �  �  �      �  Q        ����                                                                                                                                                                                                                                                                                                                           I          Q           V        Z!Vx     �  Q  [  S    �  Q  R  S    5�_�  �  �          �  T       ����                                                                                                                                                                                                                                                                                                                           I          Q           V        Z!V}   A �  S  U  \              inf.out_valid <= 1'b0;5�_�  �  �          �  T       ����                                                                                                                                                                                                                                                                                                                                                             Z!W�     �  S  U  \              inf.<= 1'b0;5�_�  �  �          �  T       ����                                                                                                                                                                                                                                                                                                                                                             Z!W�     �  S  U  \              inf.flavor_out<= 1'b0;5�_�  �  �          �  V   &    ����                                                                                                                                                                                                                                                                                                                           V   &      V   9          9    Z!W�     �  U  W  \      ;    else if (n_state == S_COMP_UPDATE || n_state == S_FILL)5�_�  �  �          �  W       ����                                                                                                                                                                                                                                                                                                                           V   &      V   9          9    Z!W�     �  V  X  \              inf.out_valid <= 1'b1;5�_�  �  �          �  W       ����                                                                                                                                                                                                                                                                                                                           V   &      V   9          9    Z!W�     �  V  X  \              inf.out_valid <= ;5�_�  �  �          �  W       ����                                                                                                                                                                                                                                                                                                                           V   &      V   9          9    Z!W�     �  V  X  \              inf.out_valid <= ();5�_�  �  �          �  W       ����                                                                                                                                                                                                                                                                                                                           V   &      V   9          9    Z!W�     �  V  X  \              inf.out_valid <= ();5�_�  �  �          �  U       ����                                                                                                                                                                                                                                                                                                                           V   &      V   9          9    Z!W�     �  T  U              end5�_�  �  �          �  S       ����                                                                                                                                                                                                                                                                                                                           U   &      U   9          9    Z!W�     �  R  T  [          if(!inf.rst_n)begin5�_�  �  �          �  L       ����                                                                                                                                                                                                                                                                                                                           U   &      U   9          9    Z!W�     �  K  L              end5�_�  �  �          �  J       ����                                                                                                                                                                                                                                                                                                                           T   &      T   9          9    Z!W�     �  I  K  Z          if(!inf.rst_n)begin5�_�  �  �          �  S       ����                                                                                                                                                                                                                                                                                                                           T   &      T   9          9    Z!W�     �  R  T  Z      #        inf.flavor_out<= no_coffee;5�_�  �  �          �  U       ����                                                                                                                                                                                                                                                                                                                           T   &      T   9          9    Z!X     �  T  V  Z      +        inf.out_valid <= () ? no_coffee : ;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                           T   &      T   9          9    Z!XO     �         [       �         Z    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                           U   &      U   9          9    Z!X`     �         [      logic not_enough = 5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                           U   &      U   9          9    Z!X`     �         [      logic not_enough = ()5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                           U   &      U   9          9    Z!Xa     �      #  [      logic not_enough = ()5�_�  �  �          �   "   )    ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�     �   !   #  ^      )                    inf.window.froth.led)5�_�  �  �          �   "   +    ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�     �   !   #  ^      -                    inf.window.froth.led) ? :5�_�  �  �          �   "   ,    ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�     �   !   #  ^      .                    inf.window.froth.led) ?  :5�_�  �  �          �   "   -    ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�     �   !   #  ^      /                    inf.window.froth.led) ? 1 :5�_�  �  �          �   "   2    ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�   B �   !   #  ^      2                    inf.window.froth.led) ? 1'b0 :5�_�  �  �          �  Y       ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�     �  X  Z  ^      ,        inf.flavor_out <= () ? no_coffee : ;5�_�  �  �          �  Y   4    ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�   C �  X  Z  ^      6        inf.flavor_out <= (not_enough) ? no_coffee : ;5�_�  �  �          �  Z       ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�     �  Y  [  ^          else5�_�  �  �          �  Z       ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!X�     �  Y  [  ^          else if 5�_�  �  �          �  Z       ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!Y     �  Y  [  ^          else if (n_state == S_FILL)5�_�  �  �          �  [       ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!Y     �  Z  [                  inf.out_valid <= 1'b0;5�_�  �  �          �  Z        ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!Y	     �  Z  \  ^              �  Z  \  ]    5�_�  �  �          �  [   #    ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!Y     �  [  ]  _          �  [  ]  ^    5�_�  �  �          �  \       ����                                                                                                                                                                                                                                                                                                                           X   &      X   9          9    Z!Y   G �  \  ^  `              �  \  ^  _    5�_�  �  �  �      �   �        ����                                                                                                                                                                                                                                                                                                                                                             Z"�     �   �   �  `       5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z"�     �   �   �  a       �   �   �  `    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z"�     �   �   �  a      assign make_coffee = 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z"�     �   �   �  a      assign make_coffee = ()5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z"�     �   �   �  a      assign make_coffee = ()5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                             Z"�     �   �   �  a      assign make_coffee = ()5�_�  �  �  �      �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  b          �   �   �  a    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      assign make_coffee = (                �   �   �  g    5�_�  �  �          �   �   .    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .assign make_coffee = (inf.window.espresso.led 5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .                      inf.window.milk.led     5�_�  �  �          �   �   .    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .assign make_coffee = (inf.window.espresso.led,5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .                      inf.window.milk.led,    5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .                      inf.window.milk.led%    5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .                      inf.window.milk.ledk    5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .                      inf.window.milk.led&    5�_�  �  �          �   �   .    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .                      inf.window.chocolate.led5�_�  �  �          �   �   .    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      .                      inf.window.froth.led    5�_�  �  �          �   �   1    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  g      1                      inf.window.froth.led  ) ? 15�_�  �  �          �   �   ,    ����                                                                                                                                                                                                                                                                                                                            �   ,          C          C    Z"�     �   �    g      �            inf.window.espresso.monitor <= (inf.window.espresso.led  )? inf.window.espresso.monitor - espresso_req  : inf.window.espresso.monitor ;   �            inf.window.milk.monitor     <= (inf.window.milk.led      )? inf.window.milk.monitor     - milk_req      : inf.window.milk.monitor     ;   �            inf.window.chocolate.monitor<= (inf.window.chocolate.led )? inf.window.chocolate.monitor- chocolate_req : inf.window.chocolate.monitor;   �            inf.window.froth.monitor    <= (inf.window.froth.led     )? inf.window.froth.monitor    - froth_req     : inf.window.froth.monitor    ;5�_�  �  �          �   �   -    ����                                                                                                                                                                                                                                                                                                                            �   ,          ,          ,    Z"   H �   �    g      {            inf.window.milk.monitor     <= ( )? inf.window.milk.monitor     - milk_req      : inf.window.milk.monitor     ;   {            inf.window.chocolate.monitor<= ( )? inf.window.chocolate.monitor- chocolate_req : inf.window.chocolate.monitor;   {            inf.window.froth.monitor    <= ( )? inf.window.froth.monitor    - froth_req     : inf.window.froth.monitor    ;�   �   �  g      {            inf.window.espresso.monitor <= ( )? inf.window.espresso.monitor - espresso_req  : inf.window.espresso.monitor ;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             Z"4�     �        h       �        g    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             Z"5	     �        h      logic fill_flag5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             Z"5
     �        h      logic fill_flag5�_�  �  �          �   ^       ����                                                                                                                                                                                                                                                                                                                                                             Z"5     �   ^   b  i       �   ^   `  h    5�_�  �  �          �   _        ����                                                                                                                                                                                                                                                                                                                            T           Z           V        Z"5#     �   _   g  k    �   _   `  k    5�_�  �  �          �   b       ����                                                                                                                                                                                                                                                                                                                            T           Z           V        Z"5&     �   a   c  r              flavor_btn_r  <= 'b0;5�_�  �  �          �   d       ����                                                                                                                                                                                                                                                                                                                            d          d   <          <    Z"5.     �   c   e  r      E    else if(n_state == S_GENERAL_REQ || n_state == S_ESPRESSO) begin 5�_�  �  �  �      �   d       ����                                                                                                                                                                                                                                                                                                                            d          d   <          <    Z"58     �   c   e  r          else if() begin 5�_�  �  �          �   d   	    ����                                                                                                                                                                                                                                                                                                                            d   	       d                 Z"5C     �   c   e  r          else if(fill_flag) begin 5�_�  �  �          �   d   
    ����                                                                                                                                                                                                                                                                                                                            d   	       d                 Z"5E     �   c   e  r      
    else  5�_�  �  �          �   e       ����                                                                                                                                                                                                                                                                                                                            d   	       d                 Z"5G     �   d   f  r      #        flavor_btn_r <= flavor_btn;5�_�  �  �          �   e       ����                                                                                                                                                                                                                                                                                                                            d   	       d                 Z"5J   I �   d   f  r      $        pre_fill_flag <= flavor_btn;5�_�  �  �          �   f       ����                                                                                                                                                                                                                                                                                                                            d   	       d                 Z"5P     �   f   h  s          �   f   h  r    5�_�  �  �          �  F       ����                                                                                                                                                                                                                                                                                                                            d   	       d                 Z"5h     �  E  G  s                  else if(fill_flag)5�_�  �  �          �  F       ����                                                                                                                                                                                                                                                                                                                            d   	       d                 Z"5m   J �  E  G  s                  else if(!fill_flag)5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                                     Z"5�     �      s      #    else if(n_state == S_FILL)begin5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                                     Z"5�   L �      s          else if()begin5�_�  �      �      �   %        ����                                                                                                                                                                                                                                                                                                                            %           &           V        Z"X�   M �   $   %          typedef enum logic[3:0]   f        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_CUSTOM_BASE,S_COMP_UPDATE,S_FILL} FSM_state;5�_�  �          �  �   %        ����                                                                                                                                                                                                                                                                                                                            %           %           V        Z"X�     �   $   '        5�_�  �          �  �   d       ����                                                                                                                                                                                                                                                                                                                            d          d   <          <    Z"55     �   d   e  r    �   c   f  r      E    else if()n_state == S_GENERAL_REQ || n_state == S_ESPRESSO begin    #        flavor_btn_r <= flavor_btn;5�_�  �          �  �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"�     �   �   �  a    �   �   �  a      .assign make_coffee = (inf.window.espresso.led    .                      inf.window.milk.led        Ealways_ff@(posedge clkinf.window.chocolate.led or negedge rst_n)begin   /    if(!inf.rst_n)begiinf.window.froth.led    n   /            inf.window.espresso.monitor <= 'b0;5�_�  �          �  �  T       ����                                                                                                                                                                                                                                                                                                                           Y   &      Y   9          9    Z!Y   D �  T  U  `       5�_�  �  �      �  �  K        ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!U�     �  K  L  S              �  K  M  T              inf.flavor_out <= 15�_�  �  �          �  L       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!U�     �  K  M  T              inf.flavor_out <= 1'b0;5�_�  �  �          �  O       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!U�     �  O  P  T          �  O  Q  U              inf.flavor_out <= 15�_�  �  �          �  P       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V     �  O  Q  U              inf.flavor_out <= 5�_�  �  �          �  P       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V     �  O  Q  U              inf.flavor_out <= ()5�_�  �  �          �  P       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V     �  O  Q  U              inf.flavor_out <= ()5�_�  �  �          �  P       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V     �  O  Q  U      ,        inf.flavor_out <= () ? no_coffee : ;5�_�  �  �          �  P   *    ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V      �  O  Q  U      -        inf.flavor_out <= () ? no_coffee :  ;5�_�  �  �          �  N   ;    ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V)     �  M  O  U      @    else if (n_state == S_COMP_UPDATE || n_state == S_FILL)begin5�_�  �  �          �  P   ,    ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V*     �  P  Q  U              �  P  R  V          end5�_�  �  �          �  R       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V-     �  Q  S  V          else begin5�_�  �  �          �  S       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V/     �  S  T  V              �  S  U  W          end5�_�  �  �          �  S       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V2     �  S  T  W       5�_�  �  �          �  T        ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!V4     �  S  U  X      (        inf.flavor_out<= inf.flavor_out;5�_�  �  �          �  M       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!VG     �  M  N  X          �  M  O  Y          else if5�_�  �              �  N       ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!VI     �  M  O  Y          else if(n_state == S_)5�_�            �  �  H        ����                                                                                                                                                                                                                                                                                                                           H          H           V        Z!U�     �  G  K        5�_�  8  :      ;  9  U       ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!Q$     �  T  V  f      always_ff@()begin5�_�  9              :  U       ����                                                                                                                                                                                                                                                                                                                           U         U   *          *    Z!Q&     �  T  V  f      always_ff@(*)begin5�_�  �                       ����                                                                                                                                                                                                                                                                                                                              8         5       V   9    Z!L�     �      J    �      J      9                    espresso_remain   <= espresso_remain;   5                    milk_remain       <= milk_remain;5�_�  �  �      �  �   �       ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!I&     �   �     +          �   �    ,          else if5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!I(     �   �    ,          else if()5�_�  �              �          ����                                                                                                                                                                                                                                                                                                                              /         /          /    Z!I8     �   �    ,          else if()5�_�  �          �  �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z!D   2 �   �   �  &      �            espresso_remain <= (c_state == S_COMP_UPDAT_OUTPUT || espresso_led  )? espresso_remain - espresso_req  : espresso_remain ;�   �     &      �            milk_remain     <= (c_state == S_COMP_UPDAT_OUTPUT || milk_led      )? milk_remain     - milk_req      : milk_remain     ;   �            chocolate_remain<= (c_state == S_COMP_UPDAT_OUTPUT || chocolate_led )? chocolate_remain- chocolate_req : chocolate_remain;   �            froth_remain    <= (c_state == S_COMP_UPDAT_OUTPUT || froth_led     )? froth_remain    - froth_req     : froth_remain    ;5�_�  w          y  x   r       ����                                                                                                                                                                                                                                                                                                                            {          ~   +          +    Z!Cj     �   r   s  '    �   q   w  '      7                if(cuespresso_weight stomize_flag)begin   %                     milk_weight        %                     chocolate_weight   %                     froth_weight        5�_�  u          w  v   r       ����                                                                                                                                                                                                                                                                                                                            x          {   +          +    Z!Cf     �   r   s  $    �   q   w  $      7                if(customize_espresso_weight flag)begin   -                             milk_weight        -                end          chocolate_weight   -                else begin   froth_weight       $                    case(flavor_btn)5�_�  T          V  U   �   6    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!A�     �   �   �  !      \        user_define_base <= (c_state == S_CUSTOM_BASE) ? ingredient_base/ sum_weight : ingre5�_�                  �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z!>�     �   �   �            else if(n_state == S_)5�_�  �          �  �           ����                                                                                                                                                                                                                                                                                                                                                             Z!-�     �               5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                                                             Z!-d     �                5�_�  o          q  p      _    ����                                                                                                                                                                                                                                                                                                                               _          `          `    Z �     �         �      rtypedef enum logic[2:0]{S_IDLE,S_INPUT,S_ESPR,S_MILK,S_CHOCO,S_FROTH,S_CUSTO_BASE,S_COMP_UPDATE_OUTPUT} FSM_state;5�_�  G          I  H   �        ����                                                                                                                                                                                                                                                                                                                            �           �   >          >    Z �     �   �   �   �    �   �   �   �      espresso_remain > espresso_req    Lmilk_remain     > milk_req     always_ff@(posedge clk or negedge rst_n)begin   6chocolate_remain> chocolate_req    if(!inf.rst_n)begin   Bfroth_remain    > froth_req                espresso_remain <= 'b0;   #            milk_remain     <= 'b0;5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �G     �   �   �   �       5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �                 Z �%     �   �   �   �    �   �   �   �      logic [9:0] espresso_req                milk_req        S//----------chocolate_req--------- COMPARE & UPDATE & OUTPUT ----------------------   :always_ff@(pfroth_req    osedge clk or negedge rst_n)begin       if(!inf.rst_n)begin5�_�  a          c  b   �       ����                                                                                                                                                                                                                                                                                                                            �   )       �   )       V   )    Z ů     �   �   �   �    �   �   �   �                  S    _FROTH:begin5�_�   �           �   �   \       ����                                                                                                                                                                                                                                                                                                                            X          ^                 Z �8     �   [   ]        5��