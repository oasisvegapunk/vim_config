Vim�UnDo� ���J,��/��s��W?�B���Z6��7�=�   d   NormalOrder norm)           )      )  )  )    Y���   ) _�                             ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  module TCCin_p05�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  module TCCin_p0[3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  module TCCin_p0[3:0], in_p15�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   module TCCin_p0[3:0], in_p1[3:0]5�_�                       '    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  'module TCCin_p0[3:0], in_p1[3:0], in_p25�_�                       +    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  ,module TCCin_p0[3:0], in_p1[3:0], in_p2[3:0]5�_�      	                 3    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  3module TCCin_p0[3:0], in_p1[3:0], in_p2[3:0], in_p35�_�      
           	      7    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  8module TCCin_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�   	              
      =    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  =module TCCin_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0], opt5�_�   
                    A    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                  Bmodule TCCin_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0], opt[1:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 : in_p05�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 : in_p0[3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 : in_p0[3:0], in_p15�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 : in_p0[3:0], in_p1[3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 : in_p0[3:0], in_p1[3:0], in_p25�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 $: in_p0[3:0], in_p1[3:0], in_p2[3:0]5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 +: in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p35�_�                       /    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                Bmodule TCCin_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0], opt[1:0]�               Output pins�                 0: in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �               Output pins�                Bmodule TCCin_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0], opt[1:0]5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                Output pins5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 0: in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 9           in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 9           in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 9           in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 9           on_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 9           on_p0[3:0], on_p1[3:0], in_p2[3:0], in_p3[3:0]5�_�                       /    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 9           on_p0[3:0], on_p1[3:0], on_p2[3:0], in_p3[3:0]5�_�                       C    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                Cmodule TCC(in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0], opt[1:0]5�_�                       9    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 9           on_p0[3:0], on_p1[3:0], on_p2[3:0], on_p3[3:0]5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 input 5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 input []5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 input []5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                 input [3:0]5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             Y��
     �                 input 5�_�   #   %           $      
    ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                 input [1:0]5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                 input [1:0]5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                Dmodule TCC(in_p0[3:0], in_p1[3:0], in_p2[3:0], in_p3[3:0], opt[1:0],5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                ?module TCC(in_p0, in_p1[3:0], in_p2[3:0], in_p3[3:0], opt[1:0],5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                :module TCC(in_p0, in_p1, in_p2[3:0], in_p3[3:0], opt[1:0],5�_�   (   *           )      %    ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                5module TCC(in_p0, in_p1, in_p2, in_p3[3:0], opt[1:0],5�_�   )   +           *      *    ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                0module TCC(in_p0, in_p1, in_p2, in_p3, opt[1:0],5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               ;           on_p0[3:0], on_p1[3:0], on_p2[3:0], on_p3[3:0]);5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               6           on_p0, on_p1[3:0], on_p2[3:0], on_p3[3:0]);5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               1           on_p0, on_p1, on_p2[3:0], on_p3[3:0]);5�_�   -   /           .      %    ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               ,           on_p0, on_p1, on_p2, on_p3[3:0]);5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                             Y��#     �                 input [1:0] 5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                             Y��+     �                 output 5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                             Y��-     �                 output [3:0]5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                             Y��.    �                 output [3:0]5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                             Y��A     �               '           on_p0, on_p1, on_p2, on_p3);5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                             Y��E    �               '           in_p0, on_p1, on_p2, on_p3);5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                             Y��L     �               '           on_p0, on_p1, on_p2, on_p3);5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                             Y��Q     �               (           out_p0, on_p1, on_p2, on_p3);5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                             Y��V     �               )           out_p0, out_p1, on_p2, on_p3);5�_�   7   9           8      #    ����                                                                                                                                                                                                                                                                                                                                                             Y��]     �               )           out_p0, out_p1,out_p2, on_p3);5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                             Y��h     �                 %output [3:0] on_p0,on_p1,on_p2,on_p3;�               5�_�   9   ;           :      )    ����                                                                                                                                                                                                                                                                                                                                                             Y��k     �                 Boutput [3:0]out_p0, out_p1,out_p2, out_p3 on_p0,on_p1,on_p2,on_p3;5�_�   :   <           ;      )    ����                                                                                                                                                                                                                                                                                                                                                             Y��l     �                 +output [3:0]out_p0, out_p1,out_p2, out_p33;5�_�   ;   =           <      )    ����                                                                                                                                                                                                                                                                                                                                                             Y��n     �               5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                             Y��p     �               *output [3:0]out_p0, out_p1,out_p2, out_p3;5�_�   =   ?           >      	    ����                                                                                                                                                                                                                                                                                                                                                             Y��p     �               *output [3:0]out_p0, out_p1,out_p2, out_p3;5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                             Y��p     �               *output [3:0]out_p0, out_p1,out_p2, out_p3;5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                             Y��q     �               *output [3:0]out_p0, out_p1,out_p2, out_p3;5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                             Y��q    �               *output [3:0]out_p0, out_p1,out_p2, out_p3;5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                             Y��x     �      	          �             5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �      	   	      parameter NO_OP = 5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �      	   	      parameter NO_OP = ''5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �      	   	      parameter NO_OP = ''5�_�   E   G           F          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �      
   	      parameter NO_OP = 25�_�   F   H           G   	       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         
                Inverse = 25�_�   G   I           H   	       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �      
                   Inverse = 2'd1,5�_�   H   J           I   	       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   	            
          �   	          5�_�   I   K           J   
       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   	                      RETROGATE = 25�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   
                      RETROGATE_INVERSE = 25�_�   K   M           L      "    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �               SpecialAdder�                     �             5�_�   L   N           M           ����                                                                                                                                                                                                                                                                                                                                                             Y��
     �               SpecialAdder5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               module SpecialAdder5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               module SpecialAdder()5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               module SpecialAdder()5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               module SpecialAdder(in,out)5�_�   Q   S           R      	    ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               module SpecialAdder(in,out);5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                             Y��      �                �             5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                             Y��#     �                   in 5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                                             Y��#     �               	    in []5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                                             Y��$     �               	    in []5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                                                             Y��'     �                   in [3:0]5�_�   W   Y           X      	    ����                                                                                                                                                                                                                                                                                                                                                             Y��'     �                   in [3:0]5�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                                                             Y��(     �                   in [3:0]5�_�   Y   [           Z          ����                                                                                                                                                                                                                                                                                                                                                             Y��*     �                   input [3:0]5�_�   Z   \           [          ����                                                                                                                                                                                                                                                                                                                                                             Y��*     �                   input [3:0]5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                                                             Y��+     �                   input [3:0]5�_�   \   ^           ]          ����                                                                                                                                                                                                                                                                                                                                                             Y��0     �                   output 5�_�   ]   _           ^          ����                                                                                                                                                                                                                                                                                                                                                             Y��1     �                   output [3:0]5�_�   ^   `           _          ����                                                                                                                                                                                                                                                                                                                                                             Y��2    �                   output [3:0]5�_�   _   a           `           ����                                                                                                                                                                                                                                                                                                                                                             Y��:     �                5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                                                             Y��>     �               module SpecialAdder(in,out);5�_�   a   c           b          ����                                                                                                                                                                                                                                                                                                                                                             Y��?     �               module SpecialAdder(in,out);5�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                                                             Y��?     �               module SpecialAdder(in,out);5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                                                             Y��@     �               module SpecialAdder(in,out);5�_�   d   f           e          ����                                                                                                                                                                                                                                                                                                                                                             Y��J     �                   input [3:0];5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                                                             Y��N     �                   input [3:0],add;5�_�   f   h           g          ����                                                                                                                                                                                                                                                                                                                                                             Y��R     �                   output [3:0];5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                                                             Y��T    �             5�_�   h   j           i           ����                                                                                                                                                                                                                                                                                                                                                             Y��V     �                5�_�   i   k           j      	    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �               	    wire 5�_�   j   l           k      
    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   wire []5�_�   k   m           l      
    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   wire []5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   wire [3:0]5�_�   m   o           n          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   input [3:0] in, add;5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                module SpecialAdder(in,out,add);5�_�   o   q           p          ����                                                                                                                                                                                                                                                                                                                                                             Y��    �                module SpecialAdder(in,out,add);5�_�   p   r           q          ����                                                                                                                                                                                                                                                                                                                                                             Y��      �               module SpecialSub(in,out,add);5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                                                             Y��!     �               module SpecialSub(in,out,);5�_�   r   t           s          ����                                                                                                                                                                                                                                                                                                                                                             Y��#     �               module SpecialSub(in,out);5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                                                             Y��&     �               module SpecialSub(in,,out);5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                                                             Y��2     �               module SpecialSub(in,,out);5�_�   u   w           v          ����                                                                                                                                                                                                                                                                                                                                                             Y��:     �                   input [3:0] in, add;�               module SpecialSub(in,sub,out);5�_�   v   x           w          ����                                                                                                                                                                                                                                                                                                                                                             Y��?     �                   input [3:0] in, add;5�_�   w   y           x          ����                                                                                                                                                                                                                                                                                                                                                             Y��A     �                   input [3:0] sub, add;5�_�   x   z           y          ����                                                                                                                                                                                                                                                                                                                                                             Y��B     �                   input [3:0] sub, add;5�_�   y   {           z          ����                                                                                                                                                                                                                                                                                                                                                             Y��E     �                   input [3:0] sub, ;5�_�   z   |           {          ����                                                                                                                                                                                                                                                                                                                                                             Y��G    �                   input [3:0] subed, ;5�_�   {   }           |          ����                                                                                                                                                                                                                                                                                                                                                             Y��K     �                   wire [3:0] tempout;5�_�   |   ~           }          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   input [3:0] subed,sub ;5�_�   }              ~          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   input [3:0] subed,sub ;5�_�   ~   �                     ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   input [3:0] subed,sub ;5�_�      �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   input [3:0] subed,sub ;5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   input [3:0] subed,sub ;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   wire [3:0] tempout = 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                   wire [3:0] tempout = 5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��     �               $    wire [3:0] tempout = subed -sub;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   �             5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[2]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[2]?5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[2] ?5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[2]) ?5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[2]) ?5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = tempout[2]) ?5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = (tempout[2]) ?5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �                   assign out = (tempout[2]) ?5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��%     �               +    assign out = (tempout[2]) ?  : tempout;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��(     �               ,    assign out = (tempout[2]) ?   : tempout;5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                             Y��0     �               3    assign out = (tempout[2]) ? tempout  : tempout;5�_�   �   �           �      (    ����                                                                                                                                                                                                                                                                                                                                                             Y��1     �               5    assign out = (tempout[2]) ? tempout[]  : tempout;5�_�   �   �           �      (    ����                                                                                                                                                                                                                                                                                                                                                             Y��2     �               5    assign out = (tempout[2]) ? tempout[]  : tempout;5�_�   �   �           �      )    ����                                                                                                                                                                                                                                                                                                                                                             Y��4     �               8    assign out = (tempout[2]) ? tempout[1:0]  : tempout;5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                             Y��4     �               8    assign out = (tempout[2]) ? tempout[1:0]  : tempout;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��5     �               8    assign out = (tempout[2]) ? tempout[1:0]  : tempout;5�_�   �   �           �      (    ����                                                                                                                                                                                                                                                                                                                                                             Y��7     �               @    assign out = (tempout[2]) ? {tempouttempout[1:0]  : tempout;5�_�   �   �           �      )    ����                                                                                                                                                                                                                                                                                                                                                             Y��8     �               B    assign out = (tempout[2]) ? {tempout[]tempout[1:0]  : tempout;5�_�   �   �           �      +    ����                                                                                                                                                                                                                                                                                                                                                             Y��:     �               C    assign out = (tempout[2]) ? {tempout[3]tempout[1:0]  : tempout;5�_�   �   �           �      -    ����                                                                                                                                                                                                                                                                                                                                                             Y��;     �               E    assign out = (tempout[2]) ? {tempout[3], tempout[1:0]  : tempout;5�_�   �   �           �      -    ����                                                                                                                                                                                                                                                                                                                                                             Y��<     �               G    assign out = (tempout[2]) ? {tempout[3], 'btempout[1:0]  : tempout;5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                                                             Y��>     �               H    assign out = (tempout[2]) ? {tempout[3], 1'btempout[1:0]  : tempout;5�_�   �   �           �      <    ����                                                                                                                                                                                                                                                                                                                                                             Y��A     �               K    assign out = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]  : tempout;5�_�   �   �           �      >    ����                                                                                                                                                                                                                                                                                                                                                             Y��A     �               K    assign out = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]  : tempout;5�_�   �   �           �      ?    ����                                                                                                                                                                                                                                                                                                                                                             Y��C     �               K    assign out = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]  : tempout;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��E     �                    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��F     �                 5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��F     �                 5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��G   	 �                 5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��Q     �                    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��R     �                �             5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��w     �               module NormalOrder5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��x     �               module NormalOrder()5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��{     �               module NormalOrder();5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �                module NormalOrder(in, out);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "       �         !    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "      module NormalOrder(in, out);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "      module NormalOrder(in, out);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "      module NormalOrder(in[], out);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "      module NormalOrder(in[], out);5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "      
    input 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "          input []5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "          input []5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "      module NormalOrder(in, out);�         "          input [3:0]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "      module NormalOrder(in, out);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "          input [3:0] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "          input [1:0] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "          input [15:0] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         "          input [15:0] 5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #      
    wire  5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #          wire [] 5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #          wire [] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #          wire [3:0] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #          wire [3:0] in_p 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #          wire [3:0] in_p[] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #          wire [3:0] in_p[] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         #          wire [3:0] in_p[0:3] 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �         %         for 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �         %      	   for() 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��     �         %      	   for() 5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                                                             Y��"     �         %      1   for(index =0 ; index <=15 ; index = index +1) 5�_�   �   �           �      .    ����                                                                                                                                                                                                                                                                                                                                                             Y��(     �         &      0   for(index =0 ; index <=15 ; index = index +1)5�_�   �   �           �      /    ����                                                                                                                                                                                                                                                                                                                                                             Y��)     �         &      0   for(index =0 ; index <=15 ; index = index +3)5�_�   �   �           �      .    ����                                                                                                                                                                                                                                                                                                                                                             Y��*   
 �         &      0   for(index =0 ; index <=15 ; index = index +3)5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��/     �         &            assign 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��5     �         &            assign in_p5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��5     �         &            assign in_p[]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��7     �         &            assign in_p[]5�_�   �   �           �      /    ����                                                                                                                                                                                                                                                                                                                                                             Y��?    �         &      1   for(index =0 ; index <=15 ; index = index + 3)5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��D     �         &      1   for(index =0 ; index <=15 ; index = index + 4)5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��P     �         &            assign in_p[index]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��[     �         &            assign in_p[index] = in5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��[     �         &            assign in_p[index] = in[]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��]     �         &            assign in_p[index] = in[]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��^     �         &      !      assign in_p[index] = in[  ]5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                                                             Y��`     �         &      &      assign in_p[index] = in[:index ]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��b     �         &      &      assign in_p[index] = in[:index ]5�_�   �   �           �      #    ����                                                                                                                                                                                                                                                                                                                                                             Y��f     �         &      .      assign in_p[index] = in[index+4 :index ]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��g     �         &      .      assign in_p[index] = in[index+4 :index ]5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                                             Y��h     �         &      /      assign in_p[index] = in[ index+4 :index ]5�_�   �   �           �      )    ����                                                                                                                                                                                                                                                                                                                                                             Y��h     �         &      /      assign in_p[index] = in[ index+4 :index ]5�_�   �   �           �      /    ����                                                                                                                                                                                                                                                                                                                                                             Y��i     �         &      /      assign in_p[index] = in[ index+4 :index ]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��l     �         &    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��n     �         '          wire [3:0] in_p[0:3];5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��n     �         '          wire [3:0] in_p[0:3];5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��q     �         '    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y��w     �         (       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��~     �         (          output 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y��~     �         (          output []5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         (          output []5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         (          output [15:0]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         (          output [15:0]5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         (    �         (    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         )          wire [3:0] in_p[0:3];5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             Y���     �         *          �         )    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             Y���    �         +          5�_�   �   �           �   "   1    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   !   #   +      1   for(index =0 ; index <=12 ; index = index + 4)5�_�   �   �           �   #   /    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   &   ,            �   #   %   +    5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -    �   #   $   -    5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   $   %           5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      0      assign in_p[index] = in[ index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      1      assign out_p[index] = in[ index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      1      assign out_p[index] = in[ index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      2      assign out_p[index] = out[ index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      #      assign out[ index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      #      assign out[ index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      "      assign out[index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      "      assign out[index+4 :index ];5�_�   �   �           �   $   !    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      "      assign out[index+4 :index ];5�_�   �   �           �   $   '    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      (      assign out[index+4 :index ] = out;5�_�   �   �           �   $   (    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      *      assign out[index+4 :index ] = out[];5�_�   �   �           �   $   (    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      *      assign out[index+4 :index ] = out[];5�_�   �   �           �   $   .    ����                                                                                                                                                                                                                                                                                                                                                             Y���    �   #   %   -      /      assign out[index+4 :index ] = out[index];5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   "   $   -      0      assign in_p[index] = in[ index+4 :index ];5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      0      assign out[index+4 :index ] = out[index] ;5�_�   �   �           �   $   %    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      0      assign out[index+4 :index ] = out[index] ;5�_�   �   �           �   $   )    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   #   %   -      0      assign out[index+4 :index ] = out[index] ;5�_�   �   �           �   $   2    ����                                                                                                                                                                                                                                                                                                                                                             Y���    �   #   %   -      3      assign out[index+4 :index ] = out[index/4 ] ;5�_�   �              �   $   '    ����                                                                                                                                                                                                                                                                                                                                                             Y��     �   #   %   -      2      assign out[index+4 :index ] = out[index/4 ];5�_�   �                $   '    ����                                                                                                                                                                                                                                                                                                                                                             Y��    �   #   %   -      2      assign out[index+4 :index ] = out[index/4 ];5�_�                  %       ����                                                                                                                                                                                                                                                                                                                                                             Y��    �   %   '   .          �   %   '   -    5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                                             Y��     �   &   (   /      //�   &   (   .    5�_�                 '       ����                                                                                                                                                                                                                                                                                                                                                             Y��3     �   '   )   /    �   '   (   /    5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y��8    �   '   )   0          wire [3:0] in_p[0:3];5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                                             Y��D     �   %   '   0      //5�_�                 '       ����                                                                                                                                                                                                                                                                                                                                                             Y��R     �   &   '              5�_�                 '       ����                                                                                                                                                                                                                                                                                                                                                             Y��W     �   '   )   0          �   '   )   /    5�_�    	             (       ����                                                                                                                                                                                                                                                                                                                                                             Y��]     �   '   )   0          SpecialSub5�_�    
          	   (       ����                                                                                                                                                                                                                                                                                                                                                             Y��a     �   '   )   0          SpecialSub(after_sub)5�_�  	            
   (       ����                                                                                                                                                                                                                                                                                                                                                             Y��b     �   '   )   0          SpecialSub(after_sub)5�_�  
               (       ����                                                                                                                                                                                                                                                                                                                                                             Y��d     �   '   )   0          SpecialSub(after_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y��g     �   '   )   0          SpecialSub(,after_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y��h     �   '   )   0          SpecialSub(,.outafter_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y��w     �   '   )   0          SpecialSub(,.out(after_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      $    SpecialSub sub0(,.out(after_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      *    SpecialSub sub0(.subed,.out(after_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      ,    SpecialSub sub0(.subed(),.out(after_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      ,    SpecialSub sub0(.subed(),.out(after_sub)5�_�                 (   !    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      1    SpecialSub sub0(.subed(),.sub,.out(after_sub)5�_�                 (   "    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      3    SpecialSub sub0(.subed(),.sub(),.out(after_sub)5�_�                 (   &    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      3    SpecialSub sub0(.subed(),.sub(),.out(after_sub)5�_�                 (   *    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      3    SpecialSub sub0(.subed(),.sub(),.out(after_sub)5�_�                 (   3    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      3    SpecialSub sub0(.subed(),.sub(),.out(after_sub)5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      4    SpecialSub sub0(.subed(),.sub(),.out(after_sub))5�_�                 (       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      8    SpecialSub sub0(.subed(in_p),.sub(),.out(after_sub))5�_�                 (        ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      :    SpecialSub sub0(.subed(in_p[]),.sub(),.out(after_sub))5�_�                 (   %    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      :    SpecialSub sub0(.subed(in_p[]),.sub(),.out(after_sub))5�_�                 (   (    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      :    SpecialSub sub0(.subed(in_p[]),.sub(),.out(after_sub))5�_�                 (   ,    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      >    SpecialSub sub0(.subed(in_p[]),.sub(in_p),.out(after_sub))5�_�                 (   -    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      @    SpecialSub sub0(.subed(in_p[]),.sub(in_p[]),.out(after_sub))5�_�                  (   -    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      @    SpecialSub sub0(.subed(in_p[]),.sub(in_p[]),.out(after_sub))5�_�    !              (   A    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   '   )   0      A    SpecialSub sub0(.subed(in_p[]),.sub(in_p[0]),.out(after_sub))5�_�     "          !   (   A    ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   (   *   0    �   (   )   0    5�_�  !  #          "   )       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   )   +   1    �   )   *   1    5�_�  "  $          #   *       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   *   ,   2    �   *   +   2    5�_�  #  %          $   )       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   (   *   3      B    SpecialSub sub0(.subed(in_p[]),.sub(in_p[0]),.out(after_sub));5�_�  $  &          %   *       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   )   +   3      B    SpecialSub sub0(.subed(in_p[]),.sub(in_p[0]),.out(after_sub));5�_�  %  '          &   +       ����                                                                                                                                                                                                                                                                                                                                                             Y���     �   *   ,   3      B    SpecialSub sub0(.subed(in_p[]),.sub(in_p[0]),.out(after_sub));5�_�  &  (          '   (       ����                                                                                                                                                                                                                                                                                                                            (          +                 Y���     �   '   -   3      B    SpecialSub sub0(.subed(in_p[]),.sub(in_p[0]),.out(after_sub));   B    SpecialSub sub1(.subed(in_p[]),.sub(in_p[0]),.out(after_sub));   B    SpecialSub sub2(.subed(in_p[]),.sub(in_p[0]),.out(after_sub));   B    SpecialSub sub3(.subed(in_p[]),.sub(in_p[0]),.out(after_sub));    �   (   )   3    5�_�  '  )          (   (   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   '   )   3      C    SpecialSub sub0(.subed(in_p[0]),.sub(in_p[0]),.out(after_sub));5�_�  (  *          )   (   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   '   )   3      C    SpecialSub sub0(.subed(in_p[0]),.sub(in_p[0]),.out(after_sub));5�_�  )  +          *   (   A    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   (   ,   3      C    SpecialSub sub1(.subed(in_p[1]),.sub(in_p[0]),.out(after_sub));   C    SpecialSub sub2(.subed(in_p[2]),.sub(in_p[0]),.out(after_sub));   C    SpecialSub sub3(.subed(in_p[3]),.sub(in_p[0]),.out(after_sub));�   '   )   3      E    SpecialSub sub0(.subed(in_p[0]),.sub(in_p[0]),.out(after_sub[]));5�_�  *  ,          +   (   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   '   -   3      E    SpecialSub sub0(.subed(in_p[0]),.sub(in_p[0]),.out(after_sub[]));   E    SpecialSub sub1(.subed(in_p[1]),.sub(in_p[0]),.out(after_sub[]));   E    SpecialSub sub2(.subed(in_p[2]),.sub(in_p[0]),.out(after_sub[]));   E    SpecialSub sub3(.subed(in_p[3]),.sub(in_p[0]),.out(after_sub[]));    �   (   )   3    5�_�  +  -          ,   ,        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���    �   +   -   3       5�_�  ,  .          -   ,   &    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���    �   ,   .   4      // �   ,   .   3    5�_�  -  /          .   -        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   4       5�_�  .  0          /   -       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   4          assign out5�_�  /  1          0   -       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   4          assign out[]5�_�  0  2          1   -       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   4          assign out[]5�_�  1  3          2   -       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   -              assign out[15]5�_�  2  4          3   -        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   4           �   -   /   4       �   -   /   3    5�_�  3  5          4   -       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   /   3          assign out_p = 45�_�  4  6          5   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   -   /   4          always@5�_�  5  7          6   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   -   /   4          always@()5�_�  6  8          7   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   -   /   4          always@()5�_�  7  9          8   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   0   2   7          end�   -   2   4          always@(*)5�_�  8  :          9   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   .   0   8              �   .   0   7    5�_�  9  ;          :   /   
    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   .   0   8      
        if5�_�  :  <          ;   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   .   0   8              if()5�_�  ;  =          <   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   .   0   8              if()5�_�  <  >          =   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   .   0   8              if(  )5�_�  =  ?          >   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8              if(  )5�_�  >  @          ?   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8              if(after_sub  )5�_�  ?  A          @   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8              if(after_sub[]  )5�_�  @  B          A   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8              if(after_sub[]  )5�_�  A  C          B   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8              if(after_sub[3]  )5�_�  B  D          C   /   !    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8      $        if(after_sub[3]>after_sub  )5�_�  C  E          D   /   "    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8      &        if(after_sub[3]>after_sub[]  )5�_�  D  F          E   /   "    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8      &        if(after_sub[3]>after_sub[]  )5�_�  E  G          F   /   $    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   .   0   8      '        if(after_sub[3]>after_sub[2]  )5�_�  F  H          G   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��*     �   .   /          ,        if(after_sub[3]>after_sub[2] && d  )5�_�  G  I          H   /        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��+     �   .   /           5�_�  H  J          I   /        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   -   /   6          always@(*)begin�   .   0   6       5�_�  I  K          J   -       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   -   /   7          �   -   /   6    5�_�  J  L          K   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   -   /   7          reg 5�_�  K  M          L   .   	    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   -   /   7      
    reg []5�_�  L  N          M   .   	    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   -   /   7      
    reg []5�_�  M  O          N   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��!     �   .   0   8          always@(*)begin�   .   1   7          always@(*)begin�   -   /   7          reg [3:0]5�_�  N  P          O   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��2     �   .   0   9          �   .   0   8    5�_�  O  Q          P   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��:     �   .   0   9          temp1 = after_sub5�_�  P  R          Q   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��:     �   .   0   9          temp1 = after_sub[]5�_�  Q  S          R   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��;     �   .   0   9          temp1 = after_sub[]5�_�  R  T          S   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��<     �   .   0   9          temp1 = after_sub[3]5�_�  S  U          T   /   $    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��?     �   .   0   9      $    temp1 = after_sub[3] - after_sub5�_�  T  V          U   /   %    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��?     �   .   0   9      &    temp1 = after_sub[3] - after_sub[]5�_�  U  W          V   /   %    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��@     �   .   0   9      &    temp1 = after_sub[3] - after_sub[]5�_�  V  X          W   /   '    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��B     �   .   0   9      '    temp1 = after_sub[3] - after_sub[2]5�_�  W  Y          X   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��G     �   -   /   9           reg [3:0] temp1,temp3,temp3;5�_�  X  Z          Y   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��G     �   -   /   9           reg [3:0] temp1,temp3,temp3;5�_�  Y  [          Z   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��H     �   -   /   9           reg [3:0] temp1,temp3,temp3;5�_�  Z  \          [   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��H     �   -   /   9           reg [3:0] temp1,temp3,temp3;5�_�  [  ]          \   .   
    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��H     �   -   /   9           reg [3:0] temp1,temp3,temp3;5�_�  \  ^          ]   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��H     �   -   /   9           reg [3:0] temp1,temp3,temp3;5�_�  ]  _          ^   .       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��H     �   -   /   9           reg [3:0] temp1,temp3,temp3;5�_�  ^  `          _   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��S     �   .   0   9      (    temp1 = after_sub[3] - after_sub[2];5�_�  _  a          `   /       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��U     �   .   0   9      (    temp1 = after_sub[3] - after_sub[2];5�_�  `  b          a   /   
    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��X     �   /   1   9    �   /   0   9    5�_�  a  c          b   0       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��Y     �   0   2   :    �   0   1   :    5�_�  b  d          c   0       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��[     �   /   1   ;      /    assign temp1 = after_sub[3] - after_sub[2];5�_�  c  e          d   1       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��]     �   0   2   ;      /    assign temp1 = after_sub[3] - after_sub[2];5�_�  d  f          e   0       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��_     �   /   1   ;      /    assign temp2 = after_sub[3] - after_sub[2];5�_�  e  g          f   0   ,    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��a     �   /   1   ;      /    assign temp2 = after_sub[2] - after_sub[2];5�_�  f  h          g   1       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��g     �   0   2   ;      /    assign temp3 = after_sub[3] - after_sub[2];5�_�  g  i          h   1       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��m     �   0   2   ;      /    assign temp3 = after_sub[0] - after_sub[2];5�_�  h  j          i   1   ,    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��o     �   0   2   ;      /    assign temp3 = after_sub[3] - after_sub[2];5�_�  i  k          j   2       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <              �   2   4   ;    5�_�  j  l          k   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <              case5�_�  k  m          l   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <              case()5�_�  l  n          m   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <              case()5�_�  m  o          n   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <              case({})5�_�  n  p          o   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <              case({})5�_�  o  q          p   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      !        case({temp1,temp2,temp3})5�_�  p  r          q   3        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      #        case({temp1,temp2,temp3[]})5�_�  q  s          r   3        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      #        case({temp1,temp2,temp3[]})5�_�  r  t          s   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      $        case({temp1,temp2,temp3[3]})5�_�  s  u          t   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      $        case({temp1,temp2,temp3[3]})5�_�  t  v          u   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      $        case({temp1,temp2,temp3[3]})5�_�  u  w          v   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      &        case({temp1,temp2[],temp3[3]})5�_�  v  x          w   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      &        case({temp1,temp2[],temp3[3]})5�_�  w  y          x   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      '        case({temp1,temp2[3],temp3[3]})5�_�  x  z          y   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      '        case({temp1,temp2[3],temp3[3]})5�_�  y  {          z   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      '        case({temp1,temp2[3],temp3[3]})5�_�  z  |          {   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      )        case({temp1[],temp2[3],temp3[3]})5�_�  {  }          |   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      )        case({temp1[],temp2[3],temp3[3]})5�_�  |  ~          }   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      *        case({temp1[3],temp2[3],temp3[3]})5�_�  }            ~   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      *        case({temp1[3],temp2[3],temp3[3]})5�_�  ~  �             3   !    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      *        case({temp1[3],temp2[3],temp3[3]})5�_�    �          �   3   '    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   4   <      *        case({temp1[3],temp2[3],temp3[3]})5�_�  �  �          �   3   *    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   2   7   <      *        case({temp1[3],temp2[3],temp3[3]})5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   @                  �   3   5   ?    5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   @                  35�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �          @          wire [3:0] out_p[0:3];5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���    �          @          reg [3:0] out_p[0:3];5�_�  �  �          �   -       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   -              assign out_p = 4'd0;5�_�  �  �          �   ,       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   ?    5�_�  �  �          �   -        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   @      //5�_�  �  �          �   -        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ,   .   @      /5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   6   @                  3'b110:5�_�  �  �          �   5       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   4   6   A                          out_p5�_�  �  �          �   5       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   4   6   A                          out_p[]5�_�  �  �          �   5       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   4   6   A                          out_p[]5�_�  �  �          �   5       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��      �   4   6   A                          out_p[3:0]5�_�  �  �          �   5   !    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��#     �   4   6   A      !                    out_p[3:0] = 5�_�  �  �          �   5   "    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��#     �   4   6   A      #                    out_p[3:0] = {}5�_�  �  �          �   5   "    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��%     �   4   6   A      #                    out_p[3:0] = {}5�_�  �  �          �   5   #    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��&     �   4   6   A      $                    out_p[3:0] = {4}5�_�  �  �          �   5   1    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��.     �   4   6   A      2                    out_p[3:0] = {4'b0, after_sub}5�_�  �  �          �   5   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��.     �   4   6   A      4                    out_p[3:0] = {4'b0, after_sub[]}5�_�  �  �          �   5   3    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��1     �   4   6   A      4                    out_p[3:0] = {4'b0, after_sub[]}5�_�  �  �          �   5   1    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��4     �   4   6   A      2                    out_p[3:0] = {4'b0, after_sub}5�_�  �  �          �   5   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��4     �   4   6   A      4                    out_p[3:0] = {4'b0, after_sub[]}5�_�  �  �          �   5   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��5     �   4   6   A      4                    out_p[3:0] = {4'b0, after_sub[]}5�_�  �  �          �   5   4    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��6     �   4   6   A      5                    out_p[3:0] = {4'b0, after_sub[1]}5�_�  �  �          �   5   ?    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��8     �   4   6   A      @                    out_p[3:0] = {4'b0, after_sub[1], after_sub}5�_�  �  �          �   5   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��8     �   4   6   A      B                    out_p[3:0] = {4'b0, after_sub[1], after_sub[]}5�_�  �  �          �   5   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��:     �   4   6   A      B                    out_p[3:0] = {4'b0, after_sub[1], after_sub[]}5�_�  �  �          �   5   B    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��:     �   4   6   A      C                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2]}5�_�  �  �          �   5   M    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��<     �   4   6   A      N                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub}5�_�  �  �          �   5   O    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��=     �   4   6   A      Q                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[3]}5�_�  �  �          �   5   Q    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��?     �   4   6   A      Q                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[3]}5�_�  �  �          �   5       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��E     �   5   8   A    �   5   6   A    5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��X     �   3   5   C                  3'b110:5�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��b     �   5   7   C                  3'b110:5�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��d     �   5   7   C                  3'b110: //5�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��q     �   5   7   C                   3'b110: // 3 > 1 > 25�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��q     �   5   7   C                   3'b110: // 3 > 1 > 25�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��q     �   5   7   C                   3'b110: // 3 > 1 > 25�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��q     �   5   7   C                   3'b110: // 3 > 1 > 25�_�  �  �          �   7   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   6   8   C      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[3]};5�_�  �  �          �   7   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   6   8   C      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[1], after_sub[3]};5�_�  �  �          �   7   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   7   :   C    �   7   8   C    5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   7   9   E                  3'b110:5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   7   9   E                  3'b110: //25�_�  �  �          �   9   N    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   8   :   E      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[3]};5�_�  �  �          �   9   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   8   :   E      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[2]};5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   7   9   E                   3'b110: // 2 > 3 > 15�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   7   9   E                   3'b010: // 2 > 3 > 15�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   E                   3'b110: // 3 > 2 > 15�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   E                   3'b010: // 3 > 2 > 15�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   E                   3'b000: // 3 > 2 > 15�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   E                   3'b001: // 3 > 2 > 15�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   E                   3'b000: // 3 > 2 > 15�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   3   5   E                   3'b001: // 3 > 2 > 15�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   5   7   E                   3'b111: // 3 > 1 > 25�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   5   7   E                   3'b011: // 3 > 1 > 25�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   7   9   E                   3'b110: // 2 > 3 > 15�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   7   9   E                   3'b100: // 2 > 3 > 15�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   9   <   E    �   9   :   E    5�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   9   ;   G                  3'b110:5�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   9   ;   G                   3'b110: // 2 > 1 > 35�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   9   ;   G                   3'b110: // 2 > 1 > 35�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   9   ;   G                   3'b110: // 2 > 1 > 35�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   9   ;   G                   3'b110: // 2 > 1 > 35�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   9   ;   G                   3'b110: // 2 > 1 > 35�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   9   ;   G                   3'b100: // 2 > 1 > 35�_�  �  �          �   ;   N    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   :   <   G      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[3]};5�_�  �  �          �   ;   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   :   <   G      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[2]};5�_�  �  �          �   ;   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   :   <   G      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[1], after_sub[2]};5�_�  �  �          �   ;   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   ;   >   G    �   ;   <   G    5�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   ;   =   I                  3'b110:5�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��     �   ;   =   I                  3'b110: // 1 > 2 >35�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��!     �   ;   =   I                   3'b110: // 1 > 2 > 35�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��!     �   ;   =   I                   3'b110: // 1 > 2 > 35�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��!     �   ;   =   I                   3'b110: // 1 > 2 > 35�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��!     �   ;   =   I                   3'b110: // 1 > 2 > 35�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��4     �   ;   =   I                   3'b110: // 1 > 2 > 35�_�  �  �          �   =   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��I     �   <   >   I      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[3]};5�_�  �  �          �   =   N    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��M     �   <   >   I      R                    out_p[3:0] = {4'b0, after_sub[3], after_sub[2], after_sub[3]};5�_�  �  �          �   >        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��O     �   >   A   I    �   >   ?   I    5�_�  �  �          �   >        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��P     �   =   >           5�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��U     �   =   ?   J                  3'b110:5�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��Y     �   =   ?   J                  3'b110: // 1 > 3 >25�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��Z     �   =   ?   J                   3'b110: // 1 > 3 > 25�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��Z     �   =   ?   J                   3'b110: // 1 > 3 > 25�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��Z     �   =   ?   J                   3'b110: // 1 > 3 > 25�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��[     �   =   ?   J                   3'b110: // 1 > 3 > 25�_�  �  �          �   >       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��[    �   =   ?   J                   3'b110: // 1 > 3 > 25�_�  �  �          �   ?   2    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��l     �   >   @   J      R                    out_p[3:0] = {4'b0, after_sub[1], after_sub[2], after_sub[3]};5�_�  �  �          �   ?   @    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��n     �   >   @   J      R                    out_p[3:0] = {4'b0, after_sub[2], after_sub[2], after_sub[3]};5�_�  �  �          �   ?   N    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��p     �   >   @   J      R                    out_p[3:0] = {4'b0, after_sub[2], after_sub[3], after_sub[3]};5�_�  �  �          �   ?   N    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   ?   B   K                      �   ?   A   J    5�_�  �  �          �   A       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   @   B   L                          out_p5�_�  �  �          �   A       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   @   B   L                          out_p[]5�_�  �  �          �   A       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   @   B   L                          out_p[]5�_�  �  �          �   A       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   @   B   L                          out_p[3:0]5�_�  �  �          �   A   #    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���    �   @   B   L      #                    out_p[3:0] = 165�_�  �  �          �   B        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   A   B           5�_�  �  �          �   C        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   B   C           5�_�  �  �          �   C       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   B   C                  5�_�  �  �          �   E        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   D   E           5�_�  �  �          �   D        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   C   D           5�_�  �  �          �   D        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �   C   D           5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��U     �       "   F       5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��`     �       "   F      //  mapping in5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��a     �       "   F      //  mapping in[]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��e     �       "   F      //  mapping in[15:12]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��~     �       "   F      //  mapping in[15:12] = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��~     �       "   F      //  mapping in[15:12] = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in[15:12] = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in = in_p[3]5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       "   F      //  mapping in = {in_p[3]5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �       !          //  mapping in = {in_p[3]5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            '   @       *   @          @    Y���     �                     integer index;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            &   @       )   @          @    Y���     �                 7    for(index =0 ; index <=12 ; index = index + 4)begin5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �      !   C      2      assign in_p[index/4] = in[ index+4 :index ];5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �      !   C      2      assign in_p[index/4] = in[ index+4 :index ];5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �      !   C    5�_�  �  �          �   #       ����                                                                                                                                                                                                                                                                                                                            &   @       )   @          @    Y���     �   "   $   D          end5�_�  �  �          �   #       ����                                                                                                                                                                                                                                                                                                                            &   @       )   @          @    Y���     �   "   #          	    ddend5�_�  �             �   "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      4      assign out[index+4 :index ] = out_p[index/4 ];5�_�  �                "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      3     assign out[index+4 :index ] = out_p[index/4 ];5�_�                  "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      2    assign out[index+4 :index ] = out_p[index/4 ];5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      3    assign out [index+4 :index ] = out_p[index/4 ];5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      "    assign out  = out_p[index/4 ];5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      "    assign out  = out_p[index/4 ];5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      $    assign out[]  = out_p[index/4 ];5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      $    assign out[]  = out_p[index/4 ];5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      (    assign out[15:0]  = out_p[index/4 ];5�_�    	             "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      (    assign out[15:0]  = out_p[index/4 ];5�_�    
          	   "   (    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      (    assign out[15:0]  = out_p[index/4 ];5�_�  	            
   "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C          assign out[15:0]  = 5�_�  
               "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C          assign out[15:0]  = {}5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C          assign out[15:0]  = {}5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C          assign out[15:0]  = {out_p}5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      !    assign out[15:0]  = {out_p[]}5�_�               "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      !    assign out[15:0]  = {out_p[]}5�_�                 "   $    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      $    assign out[15:0]  = {out_p[3:0]}5�_�                 "        ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      #    assign out[15:0]  = {out_p[3:0]5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      #    assign out[15:0]  = {out_p[3:0]5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      #    assign out[15:0]  = {out_p[3:0]5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      "    assign out[15:0]  = out_p[3:0]5�_�                 "   !    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      "    assign out[15:0]  = out_p[3:0]5�_�                 "   "    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �       "   C      0    assign in_p[index/4] = in[ index+4 :index ];�   !   #   C      "    assign out[15:0]  = out_p[3:0]5�_�                 !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �       "   C      0    assign in_p[index/4] = in[ index+4 :index ];5�_�                 !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �       "   C      0    assign in_p[index/4] = in[ index+4 :index ];5�_�                 !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �       "   C      ,    assign in_p[3:0] = in[ index+4 :index ];5�_�                 !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �       "   C      ,    assign in_p[3:0] = in[ index+4 :index ];5�_�                 !   "    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �       "   C      ,    assign in_p[3:0] = in[ index+4 :index ];5�_�                 !   %    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �       "   C      ,    assign in_p[3:0] = in[ index+4 :index ];5�_�                 !   *    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���    �       "   C      ,    assign in_p[3:0] = in[ index+4 :index ];5�_�                  !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��     �       "   C           assign in_p[3:0] = in[0:15];5�_�    !              !        ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��     �       "   C      !    assign in_p[3:0] = in[15:12];5�_�     "          !   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��     �       "   C      "    assign in_p[3:0] = in[15:12]};5�_�  !  #          "   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��     �       "   C      "    assign in_p[3:0] = in[15:12]};5�_�  "  $          #   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��     �       "   C      "    assign in_p[3:0] = in[15:12]};5�_�  #  %          $   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��      �       "   C      "    assign in_p[3:0] = in[15:12]};5�_�  $  &          %   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��!     �       "   C      #    assign in_p[3:0] = {in[15:12]};�   !   #   C      #    assign out[15:0]  = out_p[3:0];5�_�  %  '          &   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��2     �       "   C      #    assign in_p[0:3] = {in[15:12]};5�_�  &  (          '   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��2     �       "   C      #    assign in_p[0:3] = {in[15:12]};5�_�  '  )          (   !       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��2     �       "   C      #    assign in_p[0:3] = {in[15:12]};5�_�  (  *          )   !   !    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��4     �       "   C      #    assign in_p[0:3] = {in[15:12]};5�_�  )  +          *   !   $    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��7     �       "   C      &    assign in_p[0:3] = {in[15:12],in};5�_�  *  ,          +   !   %    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��7     �       "   C      (    assign in_p[0:3] = {in[15:12],in[]};5�_�  +  -          ,   !   %    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��:     �       "   C      (    assign in_p[0:3] = {in[15:12],in[]};5�_�  ,  .          -   !   *    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��=     �       "   C      ,    assign in_p[0:3] = {in[15:12],in[11:8]};5�_�  -  /          .   !   -    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��?     �       "   C      /    assign in_p[0:3] = {in[15:12],in[11:8],in};5�_�  .  0          /   !   .    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��@     �       "   C      1    assign in_p[0:3] = {in[15:12],in[11:8],in[]};5�_�  /  1          0   !   .    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��A     �       "   C      1    assign in_p[0:3] = {in[15:12],in[11:8],in[]};5�_�  0  2          1   !   2    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��C     �       "   C      4    assign in_p[0:3] = {in[15:12],in[11:8],in[7:4]};5�_�  1  3          2   !   5    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��D     �       "   C      7    assign in_p[0:3] = {in[15:12],in[11:8],in[7:4],in};5�_�  2  4          3   !   9    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��F     �       "   C      <    assign in_p[0:3] = {in[15:12],in[11:8],in[7:4],in[3:0]};5�_�  3  5          4   "   #    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��M     �   !   #   C      #    assign out[15:0]  = out_p[3:0];5�_�  4  6          5   "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��P     �   !   #   C          assign out[15:0]  =5�_�  5  7          6   "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��P     �   !   #   C          assign out[15:0]  ={}5�_�  6  8          7   "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��R     �   !   #   C          assign out[15:0]  ={}5�_�  7  9          8   "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��X     �   !   #   C          assign out[15:0]  ={out_p}5�_�  8  :          9   "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��Y     �   !   #   C      !    assign out[15:0]  ={out_p[3]}5�_�  9  ;          :   "        ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��Z     �   !   #   C      !    assign out[15:0]  ={out_p[3]}5�_�  :  <          ;   "   &    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��^     �   !   #   C      '    assign out[15:0]  ={out_p[3],out_p}5�_�  ;  =          <   "   '    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��^     �   !   #   C      )    assign out[15:0]  ={out_p[3],out_p[]}5�_�  <  >          =   "   '    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��_     �   !   #   C      )    assign out[15:0]  ={out_p[3],out_p[]}5�_�  =  ?          >   "   )    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��`     �   !   #   C      *    assign out[15:0]  ={out_p[3],out_p[2]}5�_�  >  @          ?   "   /    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��b     �   !   #   C      0    assign out[15:0]  ={out_p[3],out_p[2],out_p}5�_�  ?  A          @   "   0    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��b     �   !   #   C      2    assign out[15:0]  ={out_p[3],out_p[2],out_p[]}5�_�  @  B          A   "   0    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��c     �   !   #   C      2    assign out[15:0]  ={out_p[3],out_p[2],out_p[]}5�_�  A  C          B   "   2    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��c     �   !   #   C      3    assign out[15:0]  ={out_p[3],out_p[2],out_p[1]}5�_�  B  D          C   "   8    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��f     �   !   #   C      9    assign out[15:0]  ={out_p[3],out_p[2],out_p[1],out_p}5�_�  C  E          D   "   9    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��f     �   !   #   C      ;    assign out[15:0]  ={out_p[3],out_p[2],out_p[1],out_p[]}5�_�  D  F          E   "   9    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��g     �   !   #   C      ;    assign out[15:0]  ={out_p[3],out_p[2],out_p[1],out_p[]}5�_�  E  G          F   "   <    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��h    �   !   #   C      <    assign out[15:0]  ={out_p[3],out_p[2],out_p[1],out_p[0]}5�_�  F  H          G   "   <    ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y��}    �   "   $   C    5�_�  G  I          H          ����                                                                                                                                                                                                                                                                                                                            &   @       )   @          @    Y���     �         E            �         D    5�_�  H  J          I          ����                                                                                                                                                                                                                                                                                                                            '   @       *   @          @    Y���     �         E      always@5�_�  I  K          J          ����                                                                                                                                                                                                                                                                                                                            '   @       *   @          @    Y���     �         E      	always@()5�_�  J  L          K          ����                                                                                                                                                                                                                                                                                                                            '   @       *   @          @    Y���     �         E      	always@()5�_�  K  M          L      
    ����                                                                                                                                                                                                                                                                                                                            '   @       *   @          @    Y��2     �         E      L    assign out = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]}  : tempout;5�_�  L  N          M   *   
    ����                                                                                                                                                                                                                                                                                                                            '   @       *   @          @    Y��3     �   )   +   E      F    SpecialSub sub3(.subed(in_p[3]),.sub(in_p[0]),.out(after_sub[3]));5�_�  M  O          N      	    ����                                                                                                                                                                                                                                                                                                                            '   @       *   @          @    Y��b     �         F            �         E    5�_�  N  P          O          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��i     �         F      wire 5�_�  O  Q          P          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��i     �         F      wire []5�_�  P  R          Q          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��k     �         F      wire []5�_�  Q  S          R          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��m     �         F      wire [15:0]5�_�  R  T          S          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��o     �         F      wire [15:0];5�_�  S  U          T          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y��x     �         F      wire [15:0] stage1;5�_�  T  V          U      
    ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �         F      
always@(*)5�_�  U  W          V          ����                                                                                                                                                                                                                                                                                                                            (   @       +   @          @    Y���     �         G      always@(*)begin    �         G          �         F    5�_�  V  X          W           ����                                                                                                                                                                                                                                                                                                                            +   @       .   @          @    Y���     �         I       5�_�  W  Y          X          ����                                                                                                                                                                                                                                                                                                                            +   @       .   @          @    Y���     �         I          case5�_�  X  Z          Y      	    ����                                                                                                                                                                                                                                                                                                                            +   @       .   @          @    Y���     �         I      
    case()5�_�  Y  [          Z      	    ����                                                                                                                                                                                                                                                                                                                            +   @       .   @          @    Y���     �         I      
    case()5�_�  Z  \          [          ����                                                                                                                                                                                                                                                                                                                            +   @       .   @          @    Y���     �         I          case(opt)5�_�  [  ]          \           ����                                                                                                                                                                                                                                                                                                                            .   @       1   @          @    Y���     �         L       5�_�  \  ^          ]          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op5�_�  ]  _          ^          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op[]5�_�  ^  `          _          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op[]5�_�  _  a          `          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      wire [15:0] after_op;�         M      always@(*)begin5�_�  `  b          a          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      wire [15:0] after_op;5�_�  a  c          b          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op = 5�_�  b  d          c          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op = {}5�_�  c  e          d          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op = {}5�_�  d  f          e          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op = {in_p}5�_�  e  g          f          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op = {in_p[]}5�_�  f  h          g          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                  after_op = {in_p[]}5�_�  g  i          h          ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M                   after_op = {in_p[0]}5�_�  h  j          i      $    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      %            after_op = {in_p[0],in_p}5�_�  i  k          j      %    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      '            after_op = {in_p[0],in_p[]}5�_�  j  l          k      %    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      '            after_op = {in_p[0],in_p[]}5�_�  k  m          l      '    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      (            after_op = {in_p[0],in_p[1]}5�_�  l  n          m      ,    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      -            after_op = {in_p[0],in_p[1],in_p}5�_�  m  o          n      -    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      /            after_op = {in_p[0],in_p[1],in_p[]}5�_�  n  p          o      -    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      /            after_op = {in_p[0],in_p[1],in_p[]}5�_�  o  q          p      /    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y���     �         M      0            after_op = {in_p[0],in_p[1],in_p[2]}5�_�  p  r          q      4    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y��     �         M      5            after_op = {in_p[0],in_p[1],in_p[2],in_p}5�_�  q  s          r      5    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y��     �         M      7            after_op = {in_p[0],in_p[1],in_p[2],in_p[]}5�_�  r  t          s      5    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y��     �         M      7            after_op = {in_p[0],in_p[1],in_p[2],in_p[]}5�_�  s  u          t      8    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y��     �         M      8            after_op = {in_p[0],in_p[1],in_p[2],in_p[3]}5�_�  t  v          u      8    ����                                                                                                                                                                                                                                                                                                                            /   @       2   @          @    Y��	     �         N              �         M    5�_�  u  w          v          ����                                                                                                                                                                                                                                                                                                                            1   @       4   @          @    Y��     �         O                  after_op = 5�_�  v  x          w          ����                                                                                                                                                                                                                                                                                                                            1   @       4   @          @    Y��     �         O                  after_op = {}5�_�  w  y          x          ����                                                                                                                                                                                                                                                                                                                            1   @       4   @          @    Y��[     �         O          endcase5�_�  x  z          y          ����                                                                                                                                                                                                                                                                                                                            1   @       4   @          @    Y��[     �         O      end5�_�  y  {          z          ����                                                                                                                                                                                                                                                                                                                            1   @       4   @          @    Y���     �         P                  �         O    5�_�  z  |          {          ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q                  after_op = 5�_�  {  }          |          ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q                  after_op = {}5�_�  |  ~          }          ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q                  after_op = {}5�_�  }            ~          ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      9            after_op = {in_p[0],in_p[1],in_p[2],in_p[3]};5�_�  ~  �                    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      8            after_op = {in_p0],in_p[1],in_p[2],in_p[3]};5�_�    �          �      "    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      7            after_op = {in_p0,in_p[1],in_p[2],in_p[3]};5�_�  �  �          �      #    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      6            after_op = {in_p0,in_p1],in_p[2],in_p[3]};5�_�  �  �          �      (    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      5            after_op = {in_p0,in_p1,in_p[2],in_p[3]};5�_�  �  �          �      )    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      4            after_op = {in_p0,in_p1,in_p2],in_p[3]};5�_�  �  �          �      .    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      3            after_op = {in_p0,in_p1,in_p2,in_p[3]};5�_�  �  �          �      /    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y���     �         Q      2            after_op = {in_p0,in_p1,in_p2,in_p3]};5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                            3   @       6   @          @    Y��,     �         R          �         Q    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            6   @       9   @          @    Y��0     �         T       5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            :   @       =   @          @    Y��9     �         X      function5�_�  �  �          �      	    ����                                                                                                                                                                                                                                                                                                                            :   @       =   @          @    Y��;     �         X      	function 5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                            :   @       =   @          @    Y��;     �         X      function []5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                            :   @       =   @          @    Y��<     �         X      function []5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            :   @       =   @          @    Y��>     �         X      function [15:0]5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            :   @       =   @          @    Y��C     �         X      function [15:0] inverse5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            :   @       =   @          @    Y��C     �         X      function [15:0] inverse()5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                            ;   @       >   @          @    Y���     �         Y      
    input 5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            ;   @       >   @          @    Y���     �         Y          input []5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            ;   @       >   @          @    Y���     �         Y          input []5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            ;   @       >   @          @    Y���     �         Y          input [3:0]5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            <   @       ?   @          @    Y���     �          Z    �         Z    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            A   @       D   @          @    Y���     �                    SpecialSub 5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         !          !    Y���     �         ^      F    SpecialSub sub0(.subed(in_p[0]),.sub(in_p[0]),.out(after_sub[0]));   F    SpecialSub sub1(.subed(in_p[1]),.sub(in_p[0]),.out(after_sub[1]));   F    SpecialSub sub2(.subed(in_p[2]),.sub(in_p[0]),.out(after_sub[2]));   F    SpecialSub sub3(.subed(in_p[3]),.sub(in_p[0]),.out(after_sub[3]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         !          !    Y���     �         ^      A    SpecialSub sub0(.subed(in),.sub(in_p[0]),.out(after_sub[0]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         !          !    Y���     �         ^      $    input [3:0] inv1,inv2,inv3,inv4;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         !          !    Y���     �         ^      $    input [3:0] inv0,inv2,inv3,inv4;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         !          !    Y���     �         ^      $    input [3:0] inv0,inv1,inv3,inv4;5�_�  �  �          �      "    ����                                                                                                                                                                                                                                                                                                                                         !          !    Y���     �         ^      $    input [3:0] inv0,inv1,inv2,inv4;5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                                                       Y��     �          ^      B    SpecialSub sub0(.subed(in1),.sub(in_p[0]),.out(after_sub[0]));   A    SpecialSub sub1(.subed(in),.sub(in_p[0]),.out(after_sub[1]));   A    SpecialSub sub2(.subed(in),.sub(in_p[0]),.out(after_sub[2]));   A    SpecialSub sub3(.subed(in),.sub(in_p[0]),.out(after_sub[3]));    �         ^    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y��     �         ^      C    SpecialSub sub0(.subed(in01),.sub(in_p[0]),.out(after_sub[0]));5�_�  �  �          �      %    ����                                                                                                                                                                                                                                                                                                                               %          +          +    Y��
     �         ^      ;    SpecialSub sub0(.subed(in0),.sub(),.out(after_sub[0]));�         ^      B    SpecialSub sub0(.subed(in0),.sub(in_p[0]),.out(after_sub[0]));   B    SpecialSub sub1(.subed(in1),.sub(in_p[0]),.out(after_sub[1]));   B    SpecialSub sub2(.subed(in2),.sub(in_p[0]),.out(after_sub[2]));   B    SpecialSub sub3(.subed(in3),.sub(in_p[0]),.out(after_sub[3]));5�_�  �  �          �      &    ����                                                                                                                                                                                                                                                                                                                               %          +          +    Y��     �         ^      <    SpecialSub sub0(.subed(in0),.sub(4),.out(after_sub[0]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               %          +          +    Y���     �                ?    SpecialSub sub0(.subed(in0),.sub(4'd2),.out(after_sub[0]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               %          +          +    Y���     �         ]      ?    SpecialSub sub1(.subed(in1),.sub(4'd2),.out(after_sub[1]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �         ]      ?    SpecialSub sub2(.subed(in2),.sub(4'd2),.out(after_sub[2]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       Y���    �         ]      ?    SpecialSub sub3(.subed(in3),.sub(4'd2),.out(after_sub[3]));5�_�  �  �          �      *    ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �         ]      @    SpecialSub sub1(.subed(inv1),.sub(4'd2),.out(after_sub[1]));5�_�  �  �          �      *    ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �         ]      @    SpecialSub sub2(.subed(inv2),.sub(4'd2),.out(after_sub[2]));5�_�  �  �          �      *    ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �         ]      @    SpecialSub sub2(.subed(inv2),.sub(inv2),.out(after_sub[2]));5�_�  �  �          �      *    ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �         ]      @    SpecialSub sub1(.subed(inv1),.sub(inv1),.out(after_sub[1]));5�_�  �  �          �      *    ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �         ]      @    SpecialSub sub3(.subed(inv3),.sub(4'd2),.out(after_sub[3]));5�_�  �  �          �      .    ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �      !   ]    �         ]    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       Y���     �      !   `      @    SpecialSub sub3(.subed(inv3),.sub(inv0),.out(after_sub[3]));�          `      @    SpecialSub sub2(.subed(inv2),.sub(inv0),.out(after_sub[2]));�         `      @    SpecialSub sub1(.subed(inv1),.sub(inv0),.out(after_sub[1]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                        Y���     �      !   `      A    SpecialSub sub_1(.subed(inv1),.sub(inv0),.out(after_sub[1]));   A    SpecialSub sub_2(.subed(inv2),.sub(inv0),.out(after_sub[2]));   A    SpecialSub sub_3(.subed(inv3),.sub(inv0),.out(after_sub[3]));5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                               &          )          )    Y���     �      "   `      =    SpecialSub sub_1(.subed(),.sub(inv0),.out(after_sub[1]));   =    SpecialSub sub_2(.subed(),.sub(inv0),.out(after_sub[2]));   =    SpecialSub sub_3(.subed(),.sub(inv0),.out(after_sub[3]));    �         `    5�_�  �  �          �      &    ����                                                                                                                                                                                                                                                                                                                               1          <          <    Y��     �      "   `      A    SpecialSub sub_1(.subed(inv0),.sub(inv0),.out(after_sub[1]));   A    SpecialSub sub_2(.subed(inv0),.sub(inv0),.out(after_sub[2]));   A    SpecialSub sub_3(.subed(inv0),.sub(inv0),.out(after_sub[3]));    �         `    5�_�  �  �          �      3    ����                                                                                                                                                                                                                                                                                                                               3           6          6    Y��     �      !   `      M    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]inv0),.out(after_sub[1]));   M    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]inv0),.out(after_sub[2]));   M    SpecialSub sub_3(.subed(inv0),.sub(after_sub[3]inv0),.out(after_sub[3]));5�_�  �  �          �      :    ����                                                                                                                                                                                                                                                                                                                               :           E          E    Y��     �      !   `      I    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out(after_sub[1]));   I    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]),.out(after_sub[2]));   I    SpecialSub sub_3(.subed(inv0),.sub(after_sub[3]),.out(after_sub[3]));5�_�  �  �          �      :    ����                                                                                                                                                                                                                                                                                                                               :           E          E    Y��     �         `      =    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out());5�_�  �  �          �      A    ����                                                                                                                                                                                                                                                                                                                               :           E          E    Y��      �         `      D    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out(inverse));5�_�  �  �          �      B    ����                                                                                                                                                                                                                                                                                                                               :           E          E    Y��      �         `      F    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out(inverse[]));5�_�  �  �          �      A    ����                                                                                                                                                                                                                                                                                                                               :           E          E    Y��!     �         `      F    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out(inverse[]));5�_�  �  �          �      ;    ����                                                                                                                                                                                                                                                                                                                               :           E          E    Y��"     �         `      F    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out(inverse[]));5�_�  �  �  �      �      9    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��2     �          `      =    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]),.out());�          `    5�_�  �  �          �       9    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��4     �      !   `      =    SpecialSub sub_3(.subed(inv0),.sub(after_sub[3]),.out());�       !   `    5�_�  �  �          �      B    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��>     �         `      F    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out(inverse[]));5�_�  �  �          �      B    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��F     �          `      F    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]),.out(inverse[]));5�_�  �  �          �       B    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��H    �      !   `      F    SpecialSub sub_3(.subed(inv0),.sub(after_sub[3]),.out(inverse[]));5�_�  �  �          �      F    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��P     �          `      I    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]),.out(inverse[7:4]));5�_�  �  �          �       F    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��Q    �      !   `      I    SpecialSub sub_3(.subed(inv0),.sub(after_sub[3]),.out(inverse[3:0]));5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��W     �       !           5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��W     �       !           5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��     �                @    SpecialSub sub1(.subed(inv1),.sub(inv0),.out(after_sub[1]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��     �                @    SpecialSub sub2(.subed(inv2),.sub(inv0),.out(after_sub[2]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��     �                @    SpecialSub sub3(.subed(inv3),.sub(inv0),.out(after_sub[3]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��     �                J    SpecialSub sub_1(.subed(inv0),.sub(after_sub[1]),.out(inverse[11:8]));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��     �                J    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]),.out(inverse[7:4] ));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��     �                J    SpecialSub sub_3(.subed(inv0),.sub(after_sub[3]),.out(inverse[3:0] ));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��7     �         X    �         X    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��@     �                %    wire [3:0] tempout = subed - sub;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��C     �         Z          �         Y    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��T     �         Z          assign after_sub5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��T     �         Z          assign after_sub[]5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��V     �         Z          assign after_sub[]5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��W     �         Z          assign after_sub[1]5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��]    �         Z      $    input [3:0] inv0,inv1,inv2,inv3;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��e     �         Z          assign after_sub[1] =5�_�  �  �          �      %    ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��m     �         Z    �         Z    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��m     �         [    �         [    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��p     �         \      &    assign after_sub[1] = inv1 - inv0;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��p     �         \      &    assign after_sub[1] = inv1 - inv0;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��t     �         \      &    assign after_sub[2] = inv1 - inv0;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y��u     �         \      &    assign after_sub[3] = inv1 - inv0;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y���     �         \      &    assign after_sub[1] = inv1 - inv0;5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \      &    assign after_sub[2] = inv2 - inv0;   &    assign after_sub[3] = inv3 - inv0;�         \      &    assign after_sub[1] = inv1 - inv0;5�_�  �  �          �      &    ����                                                                                                                                                                                                                                                                                                                               &          &          &    Y���     �         \      '    assign after_sub[2] = (inv2 - inv0;   '    assign after_sub[3] = (inv3 - inv0;�         \      '    assign after_sub[1] = (inv1 - inv0;5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \      (    assign after_sub[2] = (inv2 - inv0);   (    assign after_sub[3] = (inv3 - inv0);�         \      (    assign after_sub[1] = (inv1 - inv0);5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \          wire [3:0] after_sub[0:3];5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \          wire [4:0] after_sub[0:3];5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \      L    assign out = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]}  : tempout;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \      P    assign inverse = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]}  : tempout;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \      R    assign inverse[] = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]}  : tempout;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         \      R    assign inverse[] = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]}  : tempout;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y��     �         \      W    assign inverse[15:12] = (tempout[2]) ? {tempout[3], 1'b0, tempout[1:0]}  : tempout;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y��    �         \          assign inverse[15:12] = 5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                       Y��
     �          \    �         \    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y��
     �      !   ]    �          ]    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                       Y��
     �       "   ^    �       !   ^    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y��     �          _      !    assign inverse[15:12] = inv0;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y��     �          _      !    assign inverse[15:12] = inv0;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       Y��     �          _      !    assign inverse[11:12] = inv0;�      !   _      !    assign inverse[15:12] = inv0;�       "   _      !    assign inverse[15:12] = inv0;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                       Y��     �       "   _      !    assign inverse[15: 0] = inv0;�      !   _      !    assign inverse[15: 4] = inv0;5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                                                       Y��y     �          _      !    assign inverse[11: 8] = inv0;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                      !                 Y��}     �          _      !    assign inverse[11: 8] = inv0;5�_�  �  �          �      &    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      +    assign inverse[11: 8] = (after_subinv0;5�_�  �  �          �      ,    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      1    assign inverse[11: 8] = (after_sub[ ])? inv0;5�_�  �  �          �      -    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      3    assign inverse[11: 8] = (after_sub[ ])? {}inv0;5�_�  �  �          �      6    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      <    assign inverse[11: 8] = (after_sub[ ])? {after_sub}inv0;5�_�  �  �          �      7    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      >    assign inverse[11: 8] = (after_sub[ ])? {after_sub[]}inv0;5�_�  �  �          �      8    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      >    assign inverse[11: 8] = (after_sub[ ])? {after_sub[]}inv0;5�_�  �  �          �      9    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      @    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][]}inv0;5�_�  �  �          �      9    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      @    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][]}inv0;5�_�  �  �          �      ;    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      A    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3]}inv0;5�_�  �  �          �      <    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      B    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],}inv0;5�_�  �  �          �      ?    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      F    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],'b0'}inv0;5�_�  �  �          �      <    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      F    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],'b0'}inv0;5�_�  �  �          �      ?    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      G    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0'}inv0;5�_�  �  �          �      A    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      G    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0'}inv0;5�_�  �  �          �      K    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      Q    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub}inv0;5�_�  �             �      L    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      S    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub[]}inv0;5�_�  �                   M    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      S    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub[]}inv0;5�_�                     Q    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      X    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub[][1:0]}inv0;5�_�                    S    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �      "   _      !    assign inverse[ 7: 4] = inv0;   !    assign inverse[ 3: 0] = inv0;�          _      X    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub[][1:0]}inv0;5�_�                    '    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �          _      [    assign inverse[11: 8] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;5�_�                     '    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �      !   _      [    assign inverse[ 7: 4] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;5�_�                 !   '    ����                                                                                                                                                                                                                                                                                                                                      !                 Y���     �       "   _      [    assign inverse[ 3: 0] = (after_sub[ ])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;5�_�                    )    ����                                                                                                                                                                                                                                                                                                                               )       !   )          )    Y���     �          _      [    assign inverse[11: 8] = (after_sub[1])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;5�_�                    +    ����                                                                                                                                                                                                                                                                                                                               )       !   )          )    Y���     �      "   _      [    assign inverse[ 7: 4] = (after_sub[2])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;   [    assign inverse[ 3: 0] = (after_sub[3])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;�          _      ^    assign inverse[11: 8] = (after_sub[1][2])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;5�_�    	                9    ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y���     �      #   _      ^    assign inverse[11: 8] = (after_sub[1][2])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;   ^    assign inverse[ 7: 4] = (after_sub[2][2])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;   ^    assign inverse[ 3: 0] = (after_sub[3][2])? {after_sub[][3],1'b0, after_sub[][1:0]} : inv0;    �          _    5�_�    
          	      O    ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y���     �      #   _      _    assign inverse[11: 8] = (after_sub[1][2])? {after_sub[1][3],1'b0, after_sub[][1:0]} : inv0;   _    assign inverse[ 7: 4] = (after_sub[2][2])? {after_sub[2][3],1'b0, after_sub[][1:0]} : inv0;   _    assign inverse[ 3: 0] = (after_sub[3][2])? {after_sub[3][3],1'b0, after_sub[][1:0]} : inv0;    �          _    5�_�  	            
   "        ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��     �   !   "           5�_�  
                      ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��     �         ^                  after_op = {}5�_�                        ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��     �         ^                  after_op = inverse5�_�                        ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��     �         ^                   after_op = inverse()5�_�                        ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��     �         ^      1            after_op = {in_p0,in_p1,in_p2,in_p3};5�_�                        ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��     �         ^      1            after_op = {in_p0,in_p1,in_p2,in_p3};5�_�                        ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��     �         ^      1            after_op = {in_p0,in_p1,in_p2,in_p3};5�_�                        ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��#     �         ^                   after_op = inverse()�         ^    5�_�                    9    ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��&   ! �         ^      9            after_op = inverse({in_p0,in_p1,in_p2,in_p3})5�_�                    0    ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��-   " �         ^      0            after_op = {in_p3,in_p2,in_p1,in_p0}5�_�                    0    ����                                                                                                                                                                                                                                                                                                                               '       !   '          '    Y��2     �         `              RETROGATE_INVERSE:�         _              �         ^    5�_�                        ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��B     �         `                  after_op = 5�_�                        ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��E     �         `                  after_op = inverse5�_�                        ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��E     �         `                   after_op = inverse()5�_�                         ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��F     �         `      1            after_op = {in_p3,in_p2,in_p1,in_p0};5�_�                        ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��G     �         `      1            after_op = {in_p3,in_p2,in_p1,in_p0};5�_�                        ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��M     �         `                   after_op = inverse()�         `    5�_�                    9    ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��O   # �         `      9            after_op = inverse({in_p3,in_p2,in_p1,in_p0})5�_�                    9    ����                                                                                                                                                                                                                                                                                                                            !   '       #   '          '    Y��R     �         a              �         `    5�_�                        ����                                                                                                                                                                                                                                                                                                                            #   '       %   '          '    Y��`   $ �         b                  after_op = 165�_�                        ����                                                                                                                                                                                                                                                                                                                            #   '       %   '          '    Y��g   % �         b                  after_op = 16'bz;5�_�                          ����                                                                                                                                                                                                                                                                                                                            #   '       %   '          '    Y��j     �                 5�_�    !                     ����                                                                                                                                                                                                                                                                                                                            "   '       $   '          '    Y��m   & �         b          �         a    5�_�     "          !           ����                                                                                                                                                                                                                                                                                                                            #   '       %   '          '    Y��|     �         c       �         b    5�_�  !  #          "          ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���     �         d      NormalOrder norm5�_�  "  $          #          ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���     �         d      NormalOrder norm()5�_�  #  %          $          ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���   ' �         d      NormalOrder norm()5�_�  $  &          %          ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���     �         d      NormalOrder norm(after_op, )5�_�  %  '          &          ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���     �         d      NormalOrder norm(after_op,{} )5�_�  &  (          '          ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���     �         d      NormalOrder norm(after_op,{} )5�_�  '  )          (      8    ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���     �         d      9NormalOrder norm(after_op,{out_p0,out_p1,out_p2,out_p3} )5�_�  (              )      8    ����                                                                                                                                                                                                                                                                                                                            %   '       '   '          '    Y���   ) �         d      8NormalOrder norm(after_op,{out_p0,out_p1,out_p2,out_p3})5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                                                       Y��"     �         _          assign inverse[15:12] = ;5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                               &          &          &    Y���     �         \      .    assign after_sub[1] = inv0 -(inv1 - inv0);5�_�  �  �      �  �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y���     �         \      '    assign after_sub[1] = (inv1 - inv0;5�_�  �  �          �      #    ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y���     �         \      (    assign after_sub[1] = (inv1 - inv0);5�_�  �              �          ����                                                                                                                                                                                                                                                                                                                               :          :          :    Y���     �         \      (    assign after_sub[1] = (inv1 - inv0);5�_�  �      �  �  �      :    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��/     �          `    �          `      F    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]),.out()inverse[]);5�_�  �          �  �      :    ����                                                                                                                                                                                                                                                                                                                               :           :          :    Y��$     �      !   `      <    SpecialSub sub_2(.subed(inv0),.sub(after_sub[2]),.out();   <    SpecialSub sub_3(.subed(inv0),.sub(after_sub[3]),.out();5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                               &          )          )    Y���     �         `    �      "   `      A    SpecialSub sub_1(.subed()inv0,.sub(inv0),.out(after_sub[1]));   A    SpecialSub sub_2(.subed()inv0,.sub(inv0),.out(after_sub[2]));   A    SpecialSub sub_3(.subed()inv0,.sub(inv0),.out(after_sub[3]));    5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                                                       Y���     �         ^    �          ^      C    SpecialSub sub0(.subed(in10),.sub(in_p[0]),.out(after_sub[0]));   B    SpecialSub sub1(.subed(in)1,.sub(in_p[0]),.out(after_sub[1]));   B    SpecialSub sub2(.subed(in)2,.sub(in_p[0]),.out(after_sub[2]));   B    SpecialSub sub3(.subed(in)3,.sub(in_p[0]),.out(after_sub[3]));    5�_�                 "       ����                                                                                                                                                                                                                                                                                                                            %   @       (   @          @    Y���     �   !   #   C      8    assign out[15:0]  = {out_p[3:還是禮拜天宵夜]}5��