Vim�UnDo� �(��Ƭ�P�#��L��u	��v���)"��   5                                   Z"X�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Z"X�     �       #   2    �       !   2    5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             Z"X�    �       "   4    5�_�                    !        ����                                                                                                                                                                                                                                                                                                                                                             Z"X�     �       "   2      RR5�_�                    !        ����                                                                                                                                                                                                                                                                                                                                                             Z"X�     �   !   "   2    �   !   "   2      typedef enum logic[3:0]   f        {S_IDLE,S_GENERAL_REQ,S_ESPRESSO,S_MILK,S_CHOCO,S_CUSTOM_BASE,S_COMP_UPDATE,S_FILL} FSM_state;5�_�                     #        ����                                                                                                                                                                                                                                                                                                                                                             Z"X�    �   #   $   4       5��