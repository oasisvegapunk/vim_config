Vim�UnDo� �M�$��l�m����{�q�,��r�x7��|  U   		$finish;  '        F      F  F  F    Z"V�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Z"*�     �         �      //   Module Name : PATTERN   4//   Release version : v1.0 (Release Date: May-2017)5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z"*�     �         �      O//   Module Name : PATTERN //   Release version : v1.0 (Release Date: May-2017)   //5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             Z"+�     �      �   �    �         �    5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �       	   task YOU_PASS_task;begin   U    $display ("-------------------------------------------------------------------");   U    $display ("                         Congratulations!                          ");   U    $display ("                  You have passed all patterns!                    ");   d    $display ("                 Your execution cycles = %5d cycles                ", total_latency);   p    $display ("                    Your total latency = %.1f ns                   ", total_latency*`CYCLE_TIME);   Y    $display ("-------------------------------------------------------------------");           $finish;   end endtask 5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �          task powerleakage;begin   +    if(outvalid === 1'b0 && image_out)begin   Y                $display("************************************************************");   Y                $display("*                    Power Leackage !                      *");   Y                $display("************************************************************");                   $finish;       end   end endtask5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �          	endmodule5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�      	              �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�      
           	   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�   	              
   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�   
                 �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   �   �           5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�    �   �   �           5�_�                    !        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   !   #      5�_�                    (        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   (   *      5�_�                    )        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�     �   (   )           5�_�                    (        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z"+�    �   '   (           5�_�                    /       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z",    �   /   1      5�_�                    6        ����                                                                                                                                                                                                                                                                                                                            6           9           V        Z",!     �   5   6          >// --------------  output powerleakage check -----------------   initial begin   (    forever @(negedge clk) powerleakage;   end5�_�                    5        ����                                                                                                                                                                                                                                                                                                                            6           6           V        Z",!     �   5   8        //�   5   7      5�_�                    H       ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",C     �   H   J      5�_�                    I        ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",D     �   H   I           5�_�                    O       ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",O     �   O   Q      5�_�                    P        ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",Q     �   P   R      5�_�                    Q        ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",R    �   P   Q           5�_�                    S        ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",^    �   R   T            YOU_PASS_task;5�_�                    I       ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",�     �   H   I              reset_signal_task;5�_�      !               H        ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",�     �   H   J            �   H   J      5�_�       "           !   G       ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",�     �   F   G              force clk = 0;5�_�   !   *           "   H       ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z"-     �   G   I            // Check By Yourself !!!5�_�   "   +   #       *   g       ����                                                                                                                                                                                                                                                                                                                            f          h          V       Z"-�     �   f   g          ?	for(input_idx=0;input_idx < 100 ;input_idx=input_idx+1) begin	5�_�   *   ,           +   f       ����                                                                                                                                                                                                                                                                                                                            f          g          V       Z"-�     �   e   f          	invalid = 1;5�_�   +   -           ,   f        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   e   g        *		k = $fscanf(input_file,"%d",image_in);		5�_�   ,   .           -   f       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   e   g        (k = $fscanf(input_file,"%d",image_in);		5�_�   -   /           .   f        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   e   g        (k = $fscanf(input_file,"%d",image_in);		5�_�   .   0           /   h        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   g   h          	end   5�_�   /   1           0   h       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   g   h          	invalid = 0;5�_�   0   2           1   h       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   g   h          	image_in = 'bx;5�_�   1   3           2   f        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   f   h      5�_�   2   4           3   f        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   e   g        ,    k = $fscanf(input_file,"%d",image_in);		5�_�   3   5           4   f   +    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   f   h      �   f   g      5�_�   4   6           5   g   $    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   f   h        0    k = $fscanf(input_file,"%d",inf.select_i);		5�_�   5   7           6   g   )    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   g   i      �   g   h      5�_�   6   8           7   h   $    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   g   i        .    k = $fscanf(input_file,"%d",inf.supply);		5�_�   7   9           8   h   -    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   h   j      �   h   i      5�_�   8   :           9   i   $    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   h   j        2    k = $fscanf(input_file,"%d",inf.flavor_btn);		5�_�   9   ;           :   i   0    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   i   k      5�_�   :   <           ;   i       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   i   k      �   i   j      5�_�   ;   =           <   j   $    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z".     �   i   k        5    k = $fscanf(input_file,"%d",inf.required_size);		5�_�   <   >           =   j   *    ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"..     �   j   l      5�_�   =   ?           >   k        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1;     �   j   k           5�_�   >   @           ?   k        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1;     �   j   k           5�_�   ?   A           @   k        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1G     �   j   k           5�_�   @   B           A   k       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1H     �   k   m            �   k   m      5�_�   A   C           B   l       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1J     �   k   m            if5�_�   B   D           C   l       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1h     �   k   m            if(flavor_btn == 4)5�_�   C   E           D   l       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1i     �   k   n            if(flavor_btn == 4)5�_�   D   F           E   l       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"1p     �   l   o      �   l   m      5�_�   E   G           F   l        ����                                                                                                                                                                                                                                                                                                                            l          n          V       Z"1x     �   k   l              if(flavor_btn == 4)   -    k = $fscanf(input_file,"%d",inf.ratio);		       @(negedge clk);	5�_�   F   H           G   i        ����                                                                                                                                                                                                                                                                                                                            l          l          V       Z"1{     �   i   m      �   i   j      5�_�   G   I           H   j       ����                                                                                                                                                                                                                                                                                                                            j          l                 Z"1~     �   j   m        -    k = $fscanf(input_file,"%d",inf.ratio);		       @(negedge clk);	�   i   k            if(flavor_btn == 4)5�_�   H   J           I   j   
    ����                                                                                                                                                                                                                                                                                                                            j          l                 Z"1�     �   j   l                    �   j   l      5�_�   I   K           J   k       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   j   l                for 5�_�   J   L           K   k       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   j   l                for (  )5�_�   K   M           L   l       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   k   m        1        k = $fscanf(input_file,"%d",inf.ratio);		5�_�   L   N           M   m       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   l   n                @(negedge clk);	5�_�   M   O           N   k   G    ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   j   l        G        for ( input_idx =0 ; input_idx <4 ; input_idx = input_idx + 1 )5�_�   N   P           O   m       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   m   o                    �   m   o      5�_�   O   Q           P   j       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   i   k                if(flavor_btn == 4)5�_�   P   R           Q   n   
    ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   n   p                �   n   p      5�_�   Q   S           R   k       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   j   l        P            for ( input_idx =0 ; input_idx <4 ; input_idx = input_idx + 1 )begin5�_�   R   T           S   k       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   j   l        K       for ( input_idx =0 ; input_idx <4 ; input_idx = input_idx + 1 )begin5�_�   S   U           T   k       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   j   l        K       for ( input_idx =0 ; input_idx <4 ; input_idx = input_idx + 1 )begin5�_�   T   V           U   o       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�    �   o   q      5�_�   U   W           V   p        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   o   q         5�_�   V   X           W   q       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   q   s            �   q   s      5�_�   W   Y           X   q       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   p   r        -    k = $fscanf(input_file,"%d",inf.ratio);		5�_�   X   Z           Y   r       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   q   s        end5�_�   Y   [           Z   r        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   q   s        end5�_�   Z   \           [   s       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   r   s              @(negedge clk);	5�_�   [   ]           \   q        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   q   s      �   q   r      5�_�   \   ^           ]   r       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�    �   q   s            @(negedge clk);	5�_�   ]   _           ^   m       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"1�     �   m   o                    �   m   o      5�_�   ^   `           _   n       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   m   o                    inf.select_i = 5�_�   _   a           `   n       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   m   o                    inf.select_i = 'bx'5�_�   `   b           a   n       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   m   o                    inf.select_i = 'bx'5�_�   a   c           b   n       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   n   p                    �   n   p      5�_�   b   d           c   o       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   n   p                    inf.supply   = 5�_�   c   e           d   o       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   n   p                     inf.supply   = 'bx;'5�_�   d   f           e   o        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   n   p                     inf.supply   = 'bx;'5�_�   e   g           f   o       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   o   q                    �   o   q      5�_�   f   h           g   p       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   o   q                    inf.flavor_btn = 5�_�   g   i           h   p        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   o   q        !            inf.flavor_btn = 'bx'5�_�   h   j           i   p   !    ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   o   q        !            inf.flavor_btn = 'bx'5�_�   i   k           j   p        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2     �   p   r      5�_�   j   l           k   j       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2!     �   i   k            if(flavor_btn == 4)begin5�_�   k   m           l   p       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2+     �   p   r                    �   p   r      5�_�   l   n           m   q        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"20     �   p   r                     inf.required_size = 5�_�   m   o           n   q   $    ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"21     �   p   r        %            inf.required_size = 'bx;'5�_�   n   p           o   q   %    ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"22     �   p   r        %            inf.required_size = 'bx;'5�_�   o   q           p   r        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"23     �   q   r           5�_�   p   t           q   x        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"2f     �   w   x           5�_�   q   u   r       t   e        ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"<     �   e   g      5�_�   t   v           u   f        ����                                                                                                                                                                                                                                                                                                                            k          n                 Z"<$     �   e   g         5�_�   u   w           v   f       ����                                                                                                                                                                                                                                                                                                                            k          n                 Z"<C    �   e   f              5�_�   v   x           w   e       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"<I     �   e   g      5�_�   w   y           x   f        ����                                                                                                                                                                                                                                                                                                                            k          n                 Z"<J     �   e   f           5�_�   x   {           y   e       ����                                                                                                                                                                                                                                                                                                                            j          m                 Z"<K     �   e   g      5�_�   y   |   z       {   V        ����                                                                                                                                                                                                                                                                                                                            V          b          V       Z"<�     �   U   V          task reset_signal_task; begin        #(0.5);   rst_n=0;   	#(2.0);   0	if((outvalid !== 0)||(image_out !== 'b0)) begin   @		$display ("------------------------------------------------");   @		$display ("                  RESET VIOLATION               ");   @		$display ("Output signal should be 0 after initial RESET   ");   @		$display ("------------------------------------------------");   
		$finish;   	end   	#(10);   rst_n=1;   	#(3)   release clk;   end endtask5�_�   {   }           |   L        ����                                                                                                                                                                                                                                                                                                                            V          V          V       Z"<�     �   L   N               �   L   N      5�_�   |   ~           }   M       ����                                                                                                                                                                                                                                                                                                                            W          W          V       Z"<�     �   L   M                 5�_�   }              ~   Y        ����                                                                                                                                                                                                                                                                                                                            V          V          V       Z"=�     �   Y   [      �   Y   Z      5�_�   ~   �              Z        ����                                                                                                                                                                                                                                                                                                                            Z           Z   +          +    Z"=�     �   Y   [        0    k = $fscanf(input_file,"%d",inf.select_i);		5�_�      �           �   Z        ����                                                                                                                                                                                                                                                                                                                            Z           Z   +          +    Z"=�     �   Y   [        $    k = $fscanf(input_file,"%d",);		5�_�   �   �           �   Z   ,    ����                                                                                                                                                                                                                                                                                                                            Z           Z   +          +    Z"=�     �   Z   \            �   Z   \      5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            Z           Z   +          +    Z"=�     �   Z   \            if5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            Z           Z   +          +    Z"=�     �   Z   \            if(supply_iter ! = 0)5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            Z           Z   +          +    Z"=�     �   Z   \            if(supply_iter ! = 0)5�_�   �   �           �   \       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   \   n        .    k = $fscanf(input_file,"%d",inf.supply);		   2    k = $fscanf(input_file,"%d",inf.flavor_btn);		   5    k = $fscanf(input_file,"%d",inf.required_size);		        if(inf.flavor_btn == 4)begin   L        for ( input_idx =0 ; input_idx <4 ; input_idx = input_idx + 1 )begin   5            k = $fscanf(input_file,"%d",inf.ratio);		               @(negedge clk);	               inf.select_i = 'bx;               inf.supply   = 'bx;   !            inf.flavor_btn = 'bx;   $            inf.required_size = 'bx;           end       end       else begin   1        k = $fscanf(input_file,"%d",inf.ratio);		           @(negedge clk);	       end�   [   ]        0    k = $fscanf(input_file,"%d",inf.select_i);		5�_�   �   �           �   m       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   m   o                �   m   o      5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   Z   \            if(supply_iter ! = 0)begin5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   Z   \            if(supply_iter  = 0)begin5�_�   �   �           �   [       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   Z   \            if(supply_iter = = 0)begin5�_�   �   �           �   n       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   n   p            �   n   p      5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   n   p            else5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   o   q                �   o   q      5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                            \          m                 Z"=�     �   o   q      5�_�   �   �           �   o        ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z"=�     �   o   t      �   o   p      5�_�   �   �           �   o       ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z"=�     �   o   q                �   o   q      5�_�   �   �           �   p       ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z"=�     �   o   q            for5�_�   �   �           �   p   	    ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z"=�     �   o   q            for(  )5�_�   �   �           �   p   K    ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z">     �   o   q        M    for( input_idx = 0 ; input_idx < supply_iter ; input_idx = input_idx +1 )5�_�   �   �           �   p   M    ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z">     �   o   q        M    for( input_idx = 0 ; input_idx < supply_iter ; input_idx = input_idx +1 )5�_�   �   �           �   t   8    ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z">     �   t   v                �   t   v      5�_�   �   �           �   u       ����                                                                                                                                                                                                                                                                                                                            \          _          V       Z">     �   t   v            end5�_�   �   �           �   q       ����                                                                                                                                                                                                                                                                                                                            q          t                 Z">     �   q   u        2        k = $fscanf(input_file,"%d",inf.supply);		   6        k = $fscanf(input_file,"%d",inf.flavor_btn);		   9        k = $fscanf(input_file,"%d",inf.required_size);		�   p   r        4        k = $fscanf(input_file,"%d",inf.select_i);		5�_�   �   �           �   t        ����                                                                                                                                                                                                                                                                                                                            k          l          V       Z">"     �   t   w      �   t   u      5�_�   �   �           �   x        ����                                                                                                                                                                                                                                                                                                                            k          l          V       Z">*    �   w   x           5�_�   �   �           �   !   	    ����                                                                                                                                                                                                                                                                                                                            k          l          V       Z"Q     �   !   #         �   !   #      5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"Q     �   !   #        integer ingredient5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"Q     �   !   #        integer ingredient[]5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"Q      �   !   #        integer ingredient[]5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"Q#     �   !   #        integer ingredient[1:4]5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"Q$     �   !   #        integer ingredient[1:4]5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"Q&     �   !   #        integer ingredient[0:4]5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"Q(     �   !   #        integer ingredient[0:]5�_�   �   �           �   "   5    ����                                                                                                                                                                                                                                                                                                                            l          m          V       Z"QB     �   "   $         �   "   $      5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                            m          n          V       Z"QZ     �   !   #      5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Qb     �       !          integer ans;5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                            m          n          V       Z"Qe     �   #   %         �   #   %      5�_�   �   �           �   K        ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"R#     �   K   M      5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z"R%     �   K   L              //5�_�   �   �           �   L        ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"R&     �   L   N      5�_�   �   �           �   M        ����                                                                                                                                                                                                                                                                                                                            o          p          V       Z"R'    �   L   M           5�_�   �   �   �       �   �        ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Re     �   �   �          C        for(check_i =0 ; check_i < 72 ; check_i = check_i + 1)begin5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Rl     �   �   �        +            k = $fscanf(ans_file,"%d",ans);5�_�   �   �           �   �   %    ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Rn     �   �   �      �   �   �      5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Ro     �   �   �      �   �   �      5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Ro     �   �   �       �   �   �       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Rp     �   �   �  !    �   �   �  !    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"Rp     �   �   �  "    �   �   �  "    5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"R�     �   �   �  #      (            k = $fscanf(ans_file,"%d",);5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"R�     �   �   �  #      3            k = $fscanf(ans_file,"%d",inf.window.);5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"S     �   �   �  #      :            k = $fscanf(ans_file,"%d",inf.window.monitor);5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S     �   �   �  #      C            k = $fscanf(ans_file,"%d",inf.window.espresso.monitor);5�_�   �   �   �       �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S     �   �   �  #    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S     �   �   �  $          !    		if(ans !== image_out )begin�   �   �  $    5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S#     �   �   �  $      (            k = $fscanf(ans_file,"%d",);5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S+     �   �   �  $      (            k = $fscanf(ans_file,"%d",);5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S3     �   �   �  $      (            k = $fscanf(ans_file,"%d",);5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S<     �   �   �  $      (            k = $fscanf(ans_file,"%d",);5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"SJ     �   �   �  $      (            k = $fscanf(ans_file,"%d",);5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"SN     �   �   �  $      (            k = $fscanf(ans_file,"%d",);5�_�   �   �           �   �   -    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"SR     �   �   �  $    �   �   �  $    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"SR     �   �   �  %    �   �   �  %    5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"SU     �   �   �  &      0            k = $fscanf(ans_file,"%d",milk_led);5�_�   �   �           �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"SZ     �   �   �  &      0            k = $fscanf(ans_file,"%d",milk_led);5�_�   �   �           �   �   .    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S]     �   �   �  &    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S_     �   �   �          inf.window.espresso.monitor5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S`     �   �   �  &    �   �   �  &    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"Sb     �   �   �  '      inf.window.espresso.monitor5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"Sc     �   �   �  '      inf.window.espresso.monitor5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"Sm     �   �   �  '      +             == inf.window.espresso.monitor5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"Sx     �   �   �  '      7            expresso_rem == inf.window.espresso.monitor5�_�   �   �           �   �   8    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"Sz     �   �   �  '      8            (expresso_rem == inf.window.espresso.monitor5�_�   �   �           �   �   .    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S     �   �   �  '      0            k = $fscanf(ans_file,"%d",milk_rem);5�_�   �   �           �   �   2    ����                                                                                                                                                                                                                                                                                                                            �   2       �   2          2    Z"S�     �   �   �  '      4            k = $fscanf(ans_file,"%d",milk_rem    );�   �   �  '      4            k = $fscanf(ans_file,"%d",expresso_rem);5�_�   �   �           �   �   3    ����                                                                                                                                                                                                                                                                                                                            �   2       �   2          2    Z"S�     �   �   �  '      5            k = $fscanf(ans_file,"%d",chocolate_rem);5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                            �   2       �   2          2    Z"S�     �   �   �  '      1            k = $fscanf(ans_file,"%d",froth_rem);5�_�   �   �           �   �   2    ����                                                                                                                                                                                                                                                                                                                            �   2       �   2          2    Z"S�     �   �   �  '      4            k = $fscanf(ans_file,"%d",expresso_led);5�_�   �   �           �   �   .    ����                                                                                                                                                                                                                                                                                                                            �   2       �   2          2    Z"S�     �   �   �  '      0            k = $fscanf(ans_file,"%d",milk_led);5�_�   �   �           �   �   3    ����                                                                                                                                                                                                                                                                                                                            �   2       �   2          2    Z"S�     �   �   �  '      5            k = $fscanf(ans_file,"%d",chocolate_led);5�_�   �   �           �   �   /    ����                                                                                                                                                                                                                                                                                                                            �   2       �   2          2    Z"S�     �   �   �  '      1            k = $fscanf(ans_file,"%d",froth_led);5�_�   �   �   �       �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   3       �   &          &    Z"S�     �   �   �  (                  �   �   �  '    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �   3       �   &          &    Z"S�     �   �   �  1   	                                    �   �   �  1    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �           �                   Z"S�     �   �   �  1      milk_rem         chocolate_rem    froth_rem        expresso_led     milk_led         chocolate_led    froth_led     �   �   �  1      expresso_rem  5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �           �                   Z"S�     �   �   �                       expresso_rem  5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0                   milk_rem      5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0                   chocolate_rem                 froth_rem                     expresso_led                  milk_led                      chocolate_led                 froth_led     �   �   �  0                  () milk_rem      5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0                  () milk_rem                     () chocolate_rem                () froth_rem                    () expresso_led                 () milk_led                     () chocolate_led                () froth_led     5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0                  (chocolate_rem                (froth_rem                    (expresso_led                 (milk_led                     (chocolate_led                (froth_led     �   �   �  0                  (milk_rem      5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      )            (milk_rem     == inf.window. 5�_�   �   �           �   �   8    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      9            (expresso_rem == inf.window.espresso.monitor05�_�   �   �           �   �   4    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      4            (milk_rem     == inf.window.milk.monitor5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      )            (chocolate_rem== inf.window. 5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      )            (froth_rem    == inf.window. 5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      )            (expresso_led == inf.window. 5�_�   �   �   �       �   �   4    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      4            (expresso_led == inf.window.espresso.led5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0      )            (milk_led     == inf.window. 5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      )            (chocolate_led== inf.window. 5�_�   �   �           �   �   )    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      )            (froth_led    == inf.window. 5�_�   �   �           �   �   1    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      2            (froth_led    == inf.window.froth.led)5�_�   �   �           �   �   8    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      9            (froth_led    == inf.window.froth.led       )5�_�   �   �           �   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      6            (chocolate_led== inf.window.chocolate.led)5�_�   �   �           �   �   0    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      1            (milk_led     == inf.window.milk.led)5�_�   �   �           �   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      5            (expresso_led == inf.window.espresso.led)5�_�   �   �           �   �   5    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T     �   �   �  0      6            (froth_rem    == inf.window.froth.monitor)5�_�   �   �           �   �   8    ����                                                                                                                                                                                                                                                                                                                            �   8       �   8          8    Z"T"     �   �   �  0      9            (milk_rem     == inf.window.milk.monitor    )�   �   �  0      9            (expresso_rem == inf.window.espresso.monitor)5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T8     �   �   �  0      :            (milk_rem     == inf.window.milk.monitor     )   :            (chocolate_rem== inf.window.chocolate.monitor)   :            (froth_rem    == inf.window.froth.monitor    )   :            (expresso_led == inf.window.espresso.led     )   :            (milk_led     == inf.window.milk.led         )   :            (chocolate_led== inf.window.chocolate.led    )   :            (froth_led    == inf.window.froth.led        )�   �   �  0      :            (expresso_rem == inf.window.espresso.monitor )5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"T>     �   �   �  0      <            if(expresso_rem == inf.window.espresso.monitor )   <            if(milk_rem     == inf.window.milk.monitor     )   <            if(chocolate_rem== inf.window.chocolate.monitor)   <            if(froth_rem    == inf.window.froth.monitor    )   <            if(expresso_led == inf.window.espresso.led     )   <            if(milk_led     == inf.window.milk.led         )   <            if(chocolate_led== inf.window.chocolate.led    )   <            if(froth_led    == inf.window.froth.led        )5�_�   �   �           �   �   <    ����                                                                                                                                                                                                                                                                                                                            �   ;       �   ;          ;    Z"TF     �   �   �  0      <            if(milk_rem     != inf.window.milk.monitor     )   <            if(chocolate_rem!= inf.window.chocolate.monitor)   <            if(froth_rem    != inf.window.froth.monitor    )   <            if(expresso_led != inf.window.espresso.led     )   <            if(milk_led     != inf.window.milk.led         )   <            if(chocolate_led!= inf.window.chocolate.led    )   <            if(froth_led    != inf.window.froth.led        )�   �   �  0      <            if(expresso_rem != inf.window.espresso.monitor )5�_�   �   �           �   �   A    ����                                                                                                                                                                                                                                                                                                                            �   @       �   @          @    Z"TQ     �   �   �  0      A            if(expresso_rem != inf.window.espresso.monitor )begin5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �   @       �   @          @    Z"TT     �   �   �  1    5�_�   �   �   �       �   �       ����                                                                                                                                                                                                                                                                                                                            �   4       �   4       V   @    Z"T~     �   �   �          B				$display ("                                                ");5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z"T�     �   �   �  1    �   �   �  1    5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z"T�     �   �   �           5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �             &    Z"T�     �   �   �  7      G				$display (" No.%d Pixel                                 ",check_i);5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �             &    Z"T�     �   �   �  7      ?				$display (" No.                                 ",check_i);5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �             &    Z"T�     �   �   �  7      D				$display (" Expected: %8b                               ", ans);5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                            �          �             &    Z"T�     �   �   �  7      J				$display (" Your    : %8b                               ", image_out);5�_�   �   �           �   �   >    ����                                                                                                                                                                                                                                                                                                                            �          �             &    Z"T�     �   �   �  7      D				$display (" Expected: %8d                               ", ans);5�_�   �   �           �   �   =    ����                                                                                                                                                                                                                                                                                                                            �          �   9          9    Z"T�     �   �   �  7      J				$display (" Your    : %8d                               ", image_out);   B				$display ("------------------------------------------------");�   �   �  7    5�_�   �   �           �   �   Y    ����                                                                                                                                                                                                                                                                                                                            �          �   9          9    Z"T�     �   �   �  7      e				$display (" Your    : %8d                               ",inf.window.espresso.monitor image_out);5�_�   �              �   �   Y    ����                                                                                                                                                                                                                                                                                                                            �          �   9          9    Z"T�     �   �   �  7      d				$display (" Your    : %8d                               ",inf.window.espresso.monitorimage_out);5�_�   �                �       ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  7    �   �   �  7    5�_�                  �       ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  ?      J				$display (" No.expresso_rem                                ",check_i);5�_�                 �   >    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  ?      G				$display (" No.milk_rem                                 ",check_i);5�_�                 �   @    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  ?      J				$display (" No.expresso_rem                                ",check_i);5�_�                 �   @    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  ?      I				$display (" No.expresso_rem                                "check_i);5�_�                 �   =    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  ?      @				$display (" No.milk_rem                                 ",);5�_�                 �   >    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  ?      L				$display (" Expected: %8d                               ",expresso_rem);5�_�                 �   I    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   e    Z"T�     �   �   �  ?      [				$display (" Your    : %8d                               ",inf.window.espresso.monitor);5�_�    	             �       ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   X    Z"T�     �   �   �  ?    �   �   �  ?    5�_�    
          	   �       ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   X    Z"T�     �   �   �  G      ?				$display (" No.milk_rem                                 ");5�_�  	            
   �   >    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   X    Z"T�     �   �   �  G      H				$display (" Expected: %8d                               ",milk_rem);5�_�  
               �   I    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   X    Z"U      �   �   �  G      W				$display (" Your    : %8d                               ",inf.window.milk.monitor);5�_�               �       ����                                                                                                                                                                                                                                                                                                                            �   4       �          V   @    Z"U     �   �   �  G    �   �   �  G    5�_�                 �   I    ����                                                                                                                                                                                                                                                                                                                            �   4       �          V   @    Z"U     �   �   �  O      \				$display (" Your    : %8d                               ",inf.window.chocolate.monitor);5�_�                 �   >    ����                                                                                                                                                                                                                                                                                                                            �   4       �          V   @    Z"U     �   �   �  O      M				$display (" Expected: %8d                               ",chocolate_rem);5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �   4       �          V   @    Z"U&     �   �   �  O    5�_�               �       ����                                                                                                                                                                                                                                                                                                                            �   ;       �   @          @    Z"U�     �   �   �  P    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �   ;       �   @          @    Z"U�     �   �   �  R                      �   �   �  Q    5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �   ;       �   @          @    Z"U�     �   �   �  R    5�_�               �   7    ����                                                                                                                                                                                                                                                                                                                            �   7       �   :          :    Z"U�     �   �   �  S      A            if(expresso_led != inf.window.espresso.led     )begin       A            if(milk_led     != inf.window.milk.led         )begin                      A            if(chocolate_led!= inf.window.chocolate.led    )begin       A            if(froth_led    != inf.window.froth.led        )begin5�_�                 �   8    ����                                                                                                                                                                                                                                                                                                                            �   8       �   <          <    Z"U�     �   �   �  S      =            if(expresso_led != inf.window.espresso.led )begin       =            if(milk_led     != inf.window.milk.led     )begin                      =            if(chocolate_led!= inf.window.chocolate.led)begin       =            if(froth_led    != inf.window.froth.led    )begin5�_�                 �   7    ����                                                                                                                                                                                                                                                                                                                            �   8       �   <          <    Z"U�     �   �   �  S      8            if(expresso_led != inf.window.espresso.led )    5�_�                 �   8    ����                                                                                                                                                                                                                                                                                                                            �   8       �   <          <    Z"U�     �   �   �  R      9            if(expresso_led != inf.window.espresso.led )    8            if(milk_led     != inf.window.milk.led     )5�_�                 �   9    ����                                                                                                                                                                                                                                                                                                                            �   8       �   <          <    Z"U�     �   �   �  Q      e            if(expresso_led != inf.window.espresso.led ) if(milk_led     != inf.window.milk.led     )                   5�_�                 �   e    ����                                                                                                                                                                                                                                                                                                                            �   8       �   <          <    Z"U�     �   �   �  P      f            if(expresso_led != inf.window.espresso.led ) if(milk_led     != inf.window.milk.led     )    8            if(chocolate_led!= inf.window.chocolate.led)5�_�                 �   f    ����                                                                                                                                                                                                                                                                                                                            �   8       �   <          <    Z"U�     �   �   �  O      �            if(expresso_led != inf.window.espresso.led ) if(milk_led     != inf.window.milk.led     ) if(chocolate_led!= inf.window.chocolate.led)    5�_�                 �   �    ����                                                                                                                                                                                                                                                                                                                            �   8       �   <          <    Z"U�     �   �   �  N      �            if(expresso_led != inf.window.espresso.led ) if(milk_led     != inf.window.milk.led     ) if(chocolate_led!= inf.window.chocolate.led)    8            if(froth_led    != inf.window.froth.led    )5�_�                 �   :    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) if(milk_led     != inf.window.milk.led     ) if(chocolate_led!= inf.window.chocolate.led) if(froth_led    != inf.window.froth.led    )5�_�                  �   >    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led     != inf.window.milk.led     ) if(chocolate_led!= inf.window.chocolate.led) if(froth_led    != inf.window.froth.led    )5�_�    !              �   i    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led     != inf.window.milk.led     ) if(chocolate_led!= inf.window.chocolate.led) if(froth_led    != inf.window.froth.led    )5�_�     "          !   �   F    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led     != inf.window.milk.led     ) &&(chocolate_led!= inf.window.chocolate.led) if(froth_led    != inf.window.froth.led    )5�_�  !  #          "   �   ]    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led     ) &&(chocolate_led!= inf.window.chocolate.led) if(froth_led    != inf.window.froth.led    )5�_�  "  $          #   �   �    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led ) &&(chocolate_led!= inf.window.chocolate.led) if(froth_led    != inf.window.froth.led    )5�_�  #  %          $   �   �    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led ) &&(chocolate_led!= inf.window.chocolate.led) && (froth_led    != inf.window.froth.led    )5�_�  $  &          %   �   �    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led ) &&(chocolate_led!= inf.window.chocolate.led) && (froth_led != inf.window.froth.led    )5�_�  %  '          &   �   �    ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led ) &&(chocolate_led!= inf.window.chocolate.led) && (froth_led != inf.window.froth.led )5�_�  &  (          '   �       ����                                                                                                                                                                                                                                                                                                                            �   8       �   �          <    Z"U�     �   �   �  M      �            if(expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led ) &&(chocolate_led!= inf.window.chocolate.led) && (froth_led != inf.window.froth.led ))5�_�  '  )          (   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z"U�     �   �   �  M    �   �   �  M    5�_�  (  *          )   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z"U�     �   �   �  U          B				$display ("------------------------------------------------");5�_�  )  +          *   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z"U�     �   �   �  T      >$display ("------------------------------------------------");5�_�  *  ,          +   �   �    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z"V     �   �   �  T      �            if((expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led ) &&(chocolate_led!= inf.window.chocolate.led) && (froth_led != inf.window.froth.led ))5�_�  +  -          ,   �   �    ����                                                                                                                                                                                                                                                                                                                            �          �          V       Z"V     �   �   �  T      �            if((expresso_led != inf.window.espresso.led ) && (milk_led != inf.window.milk.led ) &&(chocolate_led!= inf.window.chocolate.led) && (froth_led != inf.window.froth.led ))begi5�_�  ,  .          -   �        ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V     �   �   �       	   !    		if(ans !== image_out )begin   B				$display ("------------------------------------------------");   G				$display ("             Wrong Answer  No.%d             ",pat_cnt);   G				$display (" No.%d Pixel                                 ",check_i);   D				$display (" Expected: %8b                               ", ans);   J				$display (" Your    : %8b                               ", image_out);   B				$display ("------------------------------------------------");   				$finish;   			    end5�_�  -  /          .   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V     �   �   �  K      ?				$display (" No.chocolate_rem                            ");5�_�  .  0          /   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V     �   �   �  K      				$display (" No.");5�_�  /  1          0   �   >    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V&     �   �   �  K      I				$display (" Expected: %8d                               ",froth_rem);5�_�  0  2          1   �   >    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V,     �   �   �  K      @				$display (" Expected: %8d                               ",);5�_�  1  3          2   �   ?    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V-     �   �   �  K      B				$display (" Expected: %8d                               ",{});5�_�  2  4          3   �   ?    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V-     �   �   �  K      B				$display (" Expected: %8d                               ",{});5�_�  3  5          4   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"VH     �   �   �  K      o				$display (" Expected: %8d                               ",{expresso_led,milk_led,chocolate_led,froth_led});5�_�  4  6          5   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"VI     �   �   �  K      o				$display (" Expected: %4d                               ",{expresso_led,milk_led,chocolate_led,froth_led});5�_�  5  7          6   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"VK     �   �   �  K      X				$display (" Your    : %8d                               ",inf.window.froth.monitor);5�_�  6  8          7   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"VL     �   �   �  K      X				$display (" Your    : %8b                               ",inf.window.froth.monitor);5�_�  7  9          8   �   O    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"VU     �   �   �  K      X				$display (" Your    : %4b                               ",inf.window.froth.monitor);5�_�  8  :          9   �   >    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V^     �   �   �  K      T				$display (" Your    : %4b                               ",inf.window.froth.led);5�_�  9  ;          :   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V`     �   �   �  L      *                    inf.window.froth.led);5�_�  :  <          ;   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"Vq     �   �   �  N                          �   �   �  M    5�_�  ;  =          <   �   -    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V|     �   �   �  N      -                    {inf.window.espresso.led 5�_�  <  >          =   �   (    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V~     �   �   �  N      (                     inf.window.milk.led5�_�  =  ?          >   �   (    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V     �   �   �  N    �   �   �  N    5�_�  >  @          ?   �        ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�     �   �   �  O      )                     inf.window.milk.led,5�_�  ?  A          @   �   )    ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�    �   �   �  O      +                     inf.window.froth.led);5�_�  @  B          A   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�     �   �   �  Q                      �   �   �  P    5�_�  A  C          B   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�     �   �   �  Q    �   �   �  Q    5�_�  B  D          C   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�     �   �   �  R    �   �   �  R    5�_�  C  E          D   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�     �   �   �  S    �   �   �  S    5�_�  D  F          E   �       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�     �   �   �  T    �   �   �  T    5�_�  E              F  '       ����                                                                                                                                                                                                                                                                                                                            �           �   	       V   �    Z"V�    �  &  (  U      		$finish;5�_�                 �   7    ����                                                                                                                                                                                                                                                                                                                            �   7       �   7          7    Z"U�     �   �   �  S      =            if(expresso_led != inf.window.espresso.led )begin5�_�                 �   ;    ����                                                                                                                                                                                                                                                                                                                            �   ;       �   @          @    Z"U�     �   �   �  P      ;            if(expresso_led != inf.window.espresso.led        ;            if(milk_led     != inf.window.milk.led            ;            if(chocolate_led!= inf.window.chocolate.led    5�_�                 �   @    ����                                                                                                                                                                                                                                                                                                                            �   A       �          V   X    Z"U     �   �   �  G    �   �   �  G      E            if(froth_rem    != inf.window.froth.monitor    )beginmilk5�_�   �           �   �   �   A    ����                                                                                                                                                                                                                                                                                                                            �   @       �   @          @    Z"T^     �   �   �  2      A            if(milk_rem     != inf.window.milk.monitor     )begin               end5�_�   �           �   �   �   3    ����                                                                                                                                                                                                                                                                                                                            �          �                 Z"S�     �   �   �  0       5�_�   �           �   �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   3       �   &          &    Z"S�     �   �   �  '    �   �   �  '   	   G            (expresso_rem == inf.windowexpresso_rem  .espresso.monitor0   /    		if(ans !== image_out )beginmilk_rem         P				$display ("------------chocolate_rem ------------------------------------");   U				$display ("            froth_rem      Wrong Answer  No.%d             ",pat_cnt);   U				$display (" No.%d Pixelexpresso_led                                   ",check_i);   R				$display (" Expected: %milk_led      8b                               ", ans);   X				$display (" Your    : %chocolate_led 8b                               ", image_out);   P				$display ("            froth_led                                         ");   B				$display ("------------------------------------------------");5�_�   �           �   �   �   &    ����                                                                                                                                                                                                                                                                                                                            �   &       �   @          @    Z"S     �   �   �  #    �   �   �  #      C            k = $fscanf(ans_file,"%d",)inf.window.espresso.monitor;   !    		if(ans !== image_out )begin5�_�   �   �   �   �   �   �        ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"R=     �   �   �        5�_�   �               �   �       ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"R>     �   �   �        5�_�   �           �   �   �        ����                                                                                                                                                                                                                                                                                                                            n          o          V       Z"R:     �   �   �        5�_�   y           {   z   V        ����                                                                                                                                                                                                                                                                                                                            V          V          V       Z"<o     �   U   c        5�_�   q   s       t   r   x        ����                                                                                                                                                                                                                                                                                                                                                             Z"2k   
 �   w   y        5�_�   r               s   {       ����                                                                                                                                                                                                                                                                                                                                                             Z":�     �   z   |        5�_�   "   $       *   #   f        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-     �   e   i        5�_�   #   %           $   e       ����                                                                                                                                                                                                                                                                                                                            g          g          V       Z"-     �   e   f         5�_�   $   &           %   f        ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-L    �   e   g        5�_�   %   '           &   f       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-Z     �   f   g            �   f   h            5�_�   &   (           '   f       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   f   g            �   f   h            inf.select_i5�_�   '   )           (   g       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   g   h         5�_�   (               )   f       ����                                                                                                                                                                                                                                                                                                                            f          f          V       Z"-�     �   f   g            �   f   h            5�_�                    Z       ����                                                                                                                                                                                                                                                                                                                            8           8           V        Z",�     �   Y   [        '	if((outvalid !== 0)||( !== 'b0)) begin5��