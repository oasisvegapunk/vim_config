Vim�UnDo� �YM��;�pQ���D�[ 	+ES��`��p��4   �   !    else if(c_state == S_OP)begin   �      t   t       t   t   t    Z�     _�                  t   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��    �   �   �   �      !    else if(c_state == S_OP)begin5�_�             t      �        ����                                                                                                                                                                                                                                                                                                                                                             Z�u     �   �   �   �       �   �   �         always@5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             Z�y     �   �   �         
always@(*)5�_�                    �   	    ����                                                                                                                                                                                                                                                                                                                                                             Z�{     �   �   �         
always@(*)5�_�                     �   
    ����                                                                                                                                                                                                                                                                                                                                                             Z�{     �   �   �         always@(*)begin5�_�      !               �       ����                                                                                                                                                                                                                                                                                                                                                             Z�|     �   �   �             �   �   �        end5�_�       "           !   �       ����                                                                                                                                                                                                                                                                                                                                                             Z�~     �   �   �            �   �   �            for5�_�   !   #           "   �       ����                                                                                                                                                                                                                                                                                                                                                             Z؀     �   �   �            for(index = 0 ; index <=4)5�_�   "   $           #   �       ����                                                                                                                                                                                                                                                                                                                                                             Z،     �   �   �            for(index = 0 ; index <=4)5�_�   #   %           $   �       ����                                                                                                                                                                                                                                                                                                                                                             Z،     �   �   �            for(index = 0 ; index <=4)5�_�   $   &           %   �       ����                                                                                                                                                                                                                                                                                                                                                             Z؍     �   �   �            for(index = 1 ; index <=4)5�_�   %   '           &   �       ����                                                                                                                                                                                                                                                                                                                                                             Z؎     �   �   �            for(index = 1 ; index <=4)5�_�   &   (           '   �       ����                                                                                                                                                                                                                                                                                                                                                             Z؏     �   �   �            for(index = 1 ; index <=4)5�_�   '   )           (   �       ����                                                                                                                                                                                                                                                                                                                                                             Z؏     �   �   �        1    for(index = 1 ; index <=4 ; index = index +1)5�_�   (   *           )   �   1    ����                                                                                                                                                                                                                                                                                                                                                             Zؔ     �   �   �        6    for(index = 1 ; index <=4 ; index = index +1)begin5�_�   )   +           *   �   5    ����                                                                                                                                                                                                                                                                                                                                                             Zؕ     �   �   �                �   �   �            end5�_�   *   ,           +   �       ����                                                                                                                                                                                                                                                                                                                                                             Zؖ     �   �   �         5�_�   +   -           ,   �       ����                                                                                                                                                                                                                                                                                                                                                             Zؠ     �   �   �                �   �   �                M_OUT_REAL_mult5�_�   ,   .           -   �       ����                                                                                                                                                                                                                                                                                                                                                             Zئ     �   �   �                M_OUT_REAL_mult[]5�_�   -   /           .   �       ����                                                                                                                                                                                                                                                                                                                                                             Zئ     �   �   �                M_OUT_REAL_mult[]5�_�   .   0           /   �       ����                                                                                                                                                                                                                                                                                                                                                             Zا     �   �   �                M_OUT_REAL_mult[index]5�_�   /   1           0   �       ����                                                                                                                                                                                                                                                                                                                                                             Zب     �   �   �        .        M_OUT_REAL_mult[index] = tmp_mult_real5�_�   0   2           1   �   .    ����                                                                                                                                                                                                                                                                                                                                                             Zح     �   �   �        0        M_OUT_REAL_mult[index] = tmp_mult_real[]5�_�   1   3           2   �   /    ����                                                                                                                                                                                                                                                                                                                                                             Zح     �   �   �        0        M_OUT_REAL_mult[index] = tmp_mult_real[]5�_�   2   4           3   �   /    ����                                                                                                                                                                                                                                                                                                                                                             Zخ     �   �   �        5        M_OUT_REAL_mult[index] = tmp_mult_real[index]5�_�   3   5           4   �   5    ����                                                                                                                                                                                                                                                                                                                                                             Zذ     �   �   �        7        M_OUT_REAL_mult[index] = tmp_mult_real[index][]5�_�   4   6           5   �   6    ����                                                                                                                                                                                                                                                                                                                                                             Zذ     �   �   �        7        M_OUT_REAL_mult[index] = tmp_mult_real[index][]5�_�   5   7           6   �   6    ����                                                                                                                                                                                                                                                                                                                                                             Zش     �   �   �        ;        M_OUT_REAL_mult[index] = tmp_mult_real[index][14:6]5�_�   6   8           7   �   ;    ����                                                                                                                                                                                                                                                                                                                                                             Zظ    �   �   �        <        M_OUT_REAL_mult[index] = tmp_mult_real[index][14:6];5�_�   7   9           8   �   ;    ����                                                                                                                                                                                                                                                                                                                                                             Zغ     �   �   �      �   �   �        <        M_OUT_REAL_mult[index] = tmp_mult_real[index][14:6];5�_�   8   :           9   �       ����                                                                                                                                                                                                                                                                                                                                                             Zؼ     �   �   �        :        M_OUT_IM_mult[index] = tmp_mult_real[index][14:6];5�_�   9   ;           :   �       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   �   �        :        M_OUT_IM_mult[index] = tmp_mult_real[index][14:6];5�_�   :   <           ;   �        ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   �   �        <        M_OUT_IM_mult[index] = tmp_mcault_real[index][14:6];5�_�   ;   =           <   �       ����                                                                                                                                                                                                                                                                                                                                                             Z��    �   �   �        8        M_OUT_IM_mult[index] = tmp_mult_im[index][14:6];5�_�   <   >           =   �        ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   �   �        5�_�   =   ?           >   �        ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   �   �        */5�_�   >   @           ?   �       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   �   �        /*5�_�   ?   A           @   �       ����                                                                                                                                                                                                                                                                                                                                                             Z��    �   �   �         �   �   �        */5�_�   @   B           A   �        ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   �   �        reg [8:0] M_OUT_REAL_mult[1:4];5�_�   A   C           B   �        ����                                                                                                                                                                                                                                                                                                                                                             Z��    �   �   �        reg [8:0] M_OUT_IM_mult[1:4];5�_�   B   D           C   y        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�(     �   y   z      �   y   z        reg [8:0] M_OUT_REAL_mult[1:4];   reg [8:0] M_OUT_IM_mult[1:4];   always@(*)begin   6    for(index = 1 ; index <=4 ; index = index +1)begin   <        M_OUT_REAL_mult[index] = tmp_mult_real[index][14:6];   8        M_OUT_IM_mult[index] = tmp_mult_im[index][14:6];       end   end5�_�   C   E           D   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�+     �   �   �        /*5�_�   D   F           E   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�-     �   �   �        Iinteger_gen_8bit  rnd8_u2r(.in(tmp_sum_real[2]),.out(M_OUT_REAL_sum[2]));5�_�   E   G           F   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�5     �   �   �         �   �   �        */5�_�   F   H           G   z        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�:     �   y   {        5�_�   G   I           H   z        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�:     �   y   {        5�_�   H   J           I   x        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�;     �   w   y        reg [8:0] M_OUT_REAL_sum[1:4];5�_�   I   K           J   y        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�>     �   x   z        reg [8:0] M_OUT_IM_sum[1:4];5�_�   J   L           K   |       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�F     �   {   }        ;        M_OUT_REAL_sum[index] = tmp_mult_real[index][14:6];5�_�   K   M           L   }       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�K     �   |   ~        8        M_OUT_IM_mult[index] = tmp_mult_im[index][14:6];5�_�   L   N           M   }       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�M     �   |   ~        7        M_OUT_IM_sum[index] = tmp_mult_im[index][14:6];5�_�   M   O           N   |       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�S     �   {   }        9        M_OUT_REAL_sum[index] =tmp_sum_real[index][14:6];�   |   ~        7        M_OUT_IM_sum[index] = tmp_mult_im[index][14:6];5�_�   N   P           O   }   )    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�W     �   |   ~        :        M_OUT_IM_sum[index] = tmp_mult_icawm[index][14:6];5�_�   O   Q           P   }   *    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�Y     �   |   ~        8        M_OUT_IM_sum[index] = tmp_mult_ica[index][14:6];5�_�   P   R           Q   }       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�[     �   |   ~        5        M_OUT_IM_sum[index] =tmp_sum_im[index][14:6];5�_�   Q   S           R   }       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�a   	 �   |   ~        7        M_OUT_IM_sum[index] =  tmp_sum_im[index][14:6];5�_�   R   T           S   |   6    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�f     �   {   }        9        M_OUT_REAL_sum[index] =tmp_sum_real[index][14:3];5�_�   S   U           T   }   4    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�g     �   |   ~        7        M_OUT_IM_sum[index] =  tmp_sum_im[index][14:3];5�_�   T   V           U   |   5    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�h     �   {   }        7        M_OUT_REAL_sum[index] =tmp_sum_real[index][:3];5�_�   U   W           V   |   3    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�     �   {   }        8        M_OUT_REAL_sum[index] =tmp_sum_real[index][7:3];5�_�   V   X           W   }   3    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Zڀ    �   |   ~        6        M_OUT_IM_sum[index] =  tmp_sum_im[index][7:3];5�_�   W   Y           X   x       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Zڸ     �   w   y        %reg signed [8:0] M_OUT_REAL_sum[1:4];5�_�   X   Z           Y   y       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Zڼ    �   x   z        #reg signed [8:0] M_OUT_IM_sum[1:4];5�_�   Y   [           Z   y       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   y   z         �   y   {        reg signed tmp_r5�_�   Z   \           [   z       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   z   {      �   z   {        reg signed tmp_r5�_�   [   ]           \   {       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   z   |        reg signed tmp_i5�_�   \   ^           ]   z       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   y   {        reg signed []tmp_r5�_�   ]   _           ^   z       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   y   {        reg signed [8:0]tmp_r�   z   |        reg signed tmp_i5�_�   ^   `           _   {       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   z   |        reg signed []tmp_i5�_�   _   a           `   {       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   z   |        reg signed [8:0]tmp_i5�_�   `   b           a   {       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   {   }        always@(*)begin�   z   |        reg signed [8:0]tmp_i;5�_�   a   c           b   z       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��    �   y   {        reg signed [8:0]tmp_r;5�_�   b   d           c   {       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�    �   {   |         5�_�   c   e           d   ~       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   ~                   �   ~   �                tmp_r = 5�_�   d   f           e          ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   ~   �                tmp_r = ``5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   ~   �                tmp_r = ``5�_�   f   h           g          ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �   ~   �                tmp_r = 5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �      �      �   ~   �        )        tmp_r = tmp_sum_real[index][7:3];5�_�   h   j           i   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��     �      �                M_OUT_REAL_sum[index] =5�_�   i   l           j   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z��    �      �        &        M_OUT_REAL_sum[index] = tmp_r;5�_�   j   m   k       l          ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�     �      �         5�_�   l   n           m   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�     �   �   �      �      �        tmp_sum_im[index][7:3];5�_�   m   o           n   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�     �      �        tmp_sum_im[index][7:3];5�_�   n   p           o   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�     �      �        '              = tmp_sum_im[index][7:3];5�_�   o   q           p   �   	    ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�      �      �        +        tmp_i     = tmp_sum_im[index][7:3];5�_�   p   r           q   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�&     �      �        '        tmp_i = tmp_sum_im[index][7:3];5�_�   q   s           r   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�a     �   �   �                M_OUT_IM_sum[index] =  5�_�   r               s   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�a    �   �   �        %        M_OUT_IM_sum[index] =  tmp_i;5�_�   j           l   k          ����                                                                                                                                                                                                                                                                                                                            �           �           V        Z�	     �      �      �   ~   �        @        tmp_r = tmp_sum_real[indtmp_sum_im[index][7:3];ex][7:3];5�_�                   z        ����                                                                                                                                                                                                                                                                                                                                                             Zת     �   y   {   �      /*5�_�                    �       ����                                                                                                                                                                                                                                                                                                                                                             Z׮    �   �   �   �       �   �   �         */5�_�                    y       ����                                                                                                                                                                                                                                                                                                                                                             Z״     �   y   z          �   y   {        always@5�_�                    z       ����                                                                                                                                                                                                                                                                                                                                                             Z׺     �   y   {        
always@(*)5�_�                    z   	    ����                                                                                                                                                                                                                                                                                                                                                             Z׽     �   y   {        
always@(*)5�_�      	              z   
    ����                                                                                                                                                                                                                                                                                                                                                             Z׽     �   y   {        always@(*)begin5�_�      
           	   z       ����                                                                                                                                                                                                                                                                                                                                                             Z׾     �   z   {            �   z   |        end5�_�   	              
   z       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   {            �   z   |            if5�_�   
                 {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            if()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            if()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            M_OUT_REAL_sum = 5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            M_OUT_REAL_sum = ()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            M_OUT_REAL_sum = ()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   y   {        always@(*)begin�   z   |            M_OUT_REAL_sum = ()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            M_OUT_REAL_sum[] = ()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            M_OUT_REAL_sum[] = ()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |            M_OUT_REAL_sum[1] = ()5�_�                    {       ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |        &    M_OUT_REAL_sum[1] = (tmp_sum_real)5�_�                    {   %    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |        (    M_OUT_REAL_sum[1] = (tmp_sum_real[])5�_�                    {   &    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �   z   |        (    M_OUT_REAL_sum[1] = (tmp_sum_real[])5�_�                    {   (    ����                                                                                                                                                                                                                                                                                                                                                             Z�     �   z   |        $    M_OUT_REAL_sum[1] = tmp_sum_real5�_�                    {   $    ����                                                                                                                                                                                                                                                                                                                                                             Z�     �   z   |        &    M_OUT_REAL_sum[1] = tmp_sum_real[]5�_�                    {   %    ����                                                                                                                                                                                                                                                                                                                                                             Z�	     �   z   |        &    M_OUT_REAL_sum[1] = tmp_sum_real[]5�_�                    {   %    ����                                                                                                                                                                                                                                                                                                                                                             Z�     �   z   |        )    M_OUT_REAL_sum[1] = tmp_sum_real[7:3]5�_�                     {   )    ����                                                                                                                                                                                                                                                                                                                                                             Z�     �   z   |        *    M_OUT_REAL_sum[1] = tmp_sum_real[7:3];5�_�                    �        ����                                                                                                                                                                                                                                                                                                                                                             Z�k     �   �   �   �       �   �   �         /*5�_�                     �       ����                                                                                                                                                                                                                                                                                                                                                             Z�t    �   �   �          �   �   �        */5��