Vim�UnDo� )�8�y��-�[5���:lMR5T*):Q�8�*�]�   $   W    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;// if multiply result mantissas MSB       3      x       x   x   x    Zȵ    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Z�     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�!     �                  module FP_Mul5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�!     �                  module FP_Mul()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�"     �                  module FP_Mul()5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             Z�,     �                  *module FP_Mul(ae, am, be, bm, ce, cm ,ovf)5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             Z�,     �                  �               5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�1     �                �             5�_�      	                 
    ����                                                                                                                                                                                                                                                                                                                                                             Z�;     �               
    input 5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             Z�;     �                   input []5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             Z�<     �                   input []5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             Z�=     �                   parameter e =3;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�>     �                   parameter e =3;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�@     �                   parameter e =3;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�J     �                   input [e-1]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�M     �                   �             5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             Z�P     �               
    input 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�R     �                   input [3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�S     �                   input [3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�a     �                   output 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�a     �                   output []5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�c     �                   output []5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�f     �                   output [e-1:0]5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                                                             Z�o     �                   �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�u     �                   output 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�w     �                   output [3:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             Z�w     �                   output [3:0]5�_�                       '    ����                                                                                                                                                                                                                                                                                                                                                             Zƅ     �                   �             5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                             ZƖ     �         	          �      	       5�_�                    
   	    ����                                                                                                                                                                                                                                                                                                                                                             Zƚ     �   	            	    wire 5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             ZƝ     �   	                wire [7:0]5�_�                     
       ����                                                                                                                                                                                                                                                                                                                                                             Zƞ     �   	                wire [7:0]5�_�      !               
   ,    ����                                                                                                                                                                                                                                                                                                                                                             ZƲ     �   
                �   
          5�_�       "           !      	    ����                                                                                                                                                                                                                                                                                                                                                             Zƶ     �   
            	    wire 5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                             ZƸ     �   
                wire [3:0]5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             ZƸ     �   
                wire [3:0]5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                             Zƾ     �                   �             5�_�   $   &           %      	    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               	    wire 5�_�   %   '           &      
    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   wire []5�_�   &   (           '      
    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   wire []5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   wire [4:0]5�_�   (   *           )      #    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   �             5�_�   )   +           *      "    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   �             5�_�   *   ,           +      	    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �               	    wire 5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   wire [1:0]5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   wire [1:0]5�_�   -   /           .      2    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   �             5�_�   .   0           /           ����                                                                                                                                                                                                                                                                                                                                                             Z��    �                   �             5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �                   �             5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �                   assign sm = pm5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �                   assign sm = pm[7]5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �                   assign sm = pm[7]5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �                   assign sm = pm[7]? pm5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �                   assign sm = pm[7]? pm[]5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                             Z�     �                   assign sm = pm[7]? pm[]5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                             Z�!     �                   assign sm = pm[7]? pm[7:4]5�_�   7   9           8      #    ����                                                                                                                                                                                                                                                                                                                                                             Z�(     �               #    assign sm = pm[7]? pm[7:4] : pm5�_�   8   :           9      $    ����                                                                                                                                                                                                                                                                                                                                                             Z�(     �               %    assign sm = pm[7]? pm[7:4] : pm[]5�_�   9   ;           :      $    ����                                                                                                                                                                                                                                                                                                                                                             Z�*     �               %    assign sm = pm[7]? pm[7:4] : pm[]5�_�   :   <           ;      (    ����                                                                                                                                                                                                                                                                                                                                                             Z�-    �               (    assign sm = pm[7]? pm[7:4] : pm[6:3]5�_�   ;   =           <      R    ����                                                                                                                                                                                                                                                                                                                                                             Z�F     �                   �             5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                             Z�M     �                   assign rnd = pm5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                                                             Z�O     �                   assign rnd = pm[7]5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                             Z�O     �                   assign rnd = pm[7]5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                             Z�R     �                   assign rnd = pm[7]? pm5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                             Z�S     �                   assign rnd = pm[7]? pm[3]5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                             Z�T     �                   assign rnd = pm[7]? pm[3]5�_�   B   D           C      "    ����                                                                                                                                                                                                                                                                                                                                                             Z�W     �               "    assign rnd = pm[7]? pm[3] : pm5�_�   C   E           D      $    ����                                                                                                                                                                                                                                                                                                                                                             Z�X     �               %    assign rnd = pm[7]? pm[3] : pm[2]5�_�   D   F           E      %    ����                                                                                                                                                                                                                                                                                                                                                             Z�Y     �               %    assign rnd = pm[7]? pm[3] : pm[2]5�_�   E   G           F      A    ����                                                                                                                                                                                                                                                                                                                                                             Z�b    �                   �             5�_�   F   H           G           ����                                                                                                                                                                                                                                                                                                                                                             Z�q     �                   �             5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                             Z�u     �                   �             5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                             Zǂ     �                   // Shift the exponential5�_�   I   K           J      )    ����                                                                                                                                                                                                                                                                                                                                                             Zǌ     �                   // �             5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                                             ZǓ     �                   assign cm = sm + rnd;5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                                             Zǔ     �                   �             5�_�   L   N           M          ����                                                                                                                                                                                                                                                                                                                                                             Zǝ     �                   assign cm = xm5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                                                             ZǠ     �                   assign cm = xm[4]5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                                                             Zǡ     �                   assign cm = xm[4]5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                                                             ZǤ     �                   assign cm = xm[4] ? xm5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                                             ZǦ     �                   assign cm = xm[4] ? xm[4:1]5�_�   Q   S           R          ����                                                                                                                                                                                                                                                                                                                                                             Zǫ     �               *    // Shift the exponential according to 5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                             ZǬ    �                   // 5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                             Zǵ     �                   assign cm = xm[4] ? xm[4:1]5�_�   T   V           U      $    ����                                                                                                                                                                                                                                                                                                                                                             ZǸ     �               $    assign cm = xm[4] ? xm[4:1] : xm5�_�   U   W           V      (    ����                                                                                                                                                                                                                                                                                                                                                             ZǺ     �               )    assign cm = xm[4] ? xm[4:1] : xm[3:0]5�_�   V   X           W      )    ����                                                                                                                                                                                                                                                                                                                                                             ZǺ    �               )    assign cm = xm[4] ? xm[4:1] : xm[3:0]5�_�   W   Y           X      )    ����                                                                                                                                                                                                                                                                                                                                                             ZǾ     �                   �             5�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !          // �              5�_�   Y   [           Z          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !          assign 5�_�   Z   \           [          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !          assign {}5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                                                             Z��    �         !          assign {}5�_�   \   ^           ]          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !          assign {oe,ce}5�_�   ]   _           ^          ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !          assign {oe,ce} = ae + be  +5�_�   ^   `           _           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !      !    assign {oe,ce} = ae + be  +()5�_�   _   a           `           ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !      !    assign {oe,ce} = ae + be  +()5�_�   `   b           a      "    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !      #    assign {oe,ce} = ae + be  +(pm)5�_�   a   c           b      $    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !      &    assign {oe,ce} = ae + be  +(pm[7])5�_�   b   d           c      %    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !      &    assign {oe,ce} = ae + be  +(pm[7])5�_�   c   e           d      *    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !      +    assign {oe,ce} = ae + be  +(pm[7] | xm)5�_�   d   f           e      ,    ����                                                                                                                                                                                                                                                                                                                                                             Z��     �         !      .    assign {oe,ce} = ae + be  +(pm[7] | xm[4])5�_�   e   g           f      .    ����                                                                                                                                                                                                                                                                                                                                                             Z��    �         !      .    assign {oe,ce} = ae + be  +(pm[7] | xm[4])5�_�   f   h           g      2    ����                                                                                                                                                                                                                                                                                                                                                             Z�     �          "          �          !    5�_�   g   i           h      3    ����                                                                                                                                                                                                                                                                                                                                                             Z�     �         "      3    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;5�_�   h   j           i      F    ����                                                                                                                                                                                                                                                                                                                                                             Z�B     �         "      F    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;// if mantissas MSB5�_�   i   k           j      B    ����                                                                                                                                                                                                                                                                                                                                                             Z�E     �         "      F    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;// if mantissas MSB5�_�   j   l           k      8    ����                                                                                                                                                                                                                                                                                                                                                             Z�F     �         "      F    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;// if mantissas MSB5�_�   k   m           l      9    ����                                                                                                                                                                                                                                                                                                                                                             Z�G     �         "      F    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;// if mantissas MSB5�_�   l   n           m      V    ����                                                                                                                                                                                                                                                                                                                                                             Z�N     �          #      8    // -1 because if MSB is zero, we shift the mantissas�          "      V    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;// if multiply result mantissas MSB5�_�   m   o           n      .    ����                                                                                                                                                                                                                                                                                                                                                             ZȆ     �          #      8    // -1 because if MSB is zero, we shift the mantissas5�_�   n   p           o      *    ����                                                                                                                                                                                                                                                                                                                                                             ZȆ     �          #      8    // -1 because if MSB is zero, we shift the mantissas5�_�   o   q           p      +    ����                                                                                                                                                                                                                                                                                                                                                             Zȉ     �          #      8    // -1 because if MSB is zero, we shift the mantissas5�_�   p   r           q      5    ����                                                                                                                                                                                                                                                                                                                                                             Zȋ     �          #      =    // -1 because if MSB is zero, we shift left the mantissas5�_�   q   s           r      7    ����                                                                                                                                                                                                                                                                                                                                                             Zȋ     �      !   #      =    // -1 because if MSB is zero, we shift left the mantissas5�_�   r   t           s           ����                                                                                                                                                                                                                                                                                                                                                             ZȖ   	 �          $      N    // -1 because if MSB is zero, we shift left the mantissas, so decrease the   exponential�      !   $              // exponential5�_�   s   u           t      N    ����                                                                                                                                                                                                                                                                                                                                                             ZȞ     �      !   #    5�_�   t   v           u       	    ����                                                                                                                                                                                                                                                                                                                                                             Zȟ     �      !   $              // 5�_�   u   w           v           ����                                                                                                                                                                                                                                                                                                                                                             ZȠ     �      !   $              // 5�_�   v   x           w           ����                                                                                                                                                                                                                                                                                                                                                             Zȡ   
 �      !   $          // 5�_�   w               x      3    ����                                                                                                                                                                                                                                                                                                                                                             Zȴ    �         $      W    assign {oe,ce} = ae + be  +(pm[7] | xm[4]) - 1;// if multiply result mantissas MSB 5��